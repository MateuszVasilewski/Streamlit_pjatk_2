��3E     �sklearn.ensemble._forest��RandomForestClassifier���)��}�(�base_estimator��sklearn.tree._classes��DecisionTreeClassifier���)��}�(�	criterion��gini��splitter��best��	max_depth�N�min_samples_split�K�min_samples_leaf�K�min_weight_fraction_leaf�G        �max_features�N�max_leaf_nodes�N�random_state�N�min_impurity_decrease�G        �class_weight�N�	ccp_alpha�G        �_sklearn_version��1.0.1�ub�n_estimators�K
�estimator_params�(hhhhhhhhhht��	bootstrap���	oob_score���n_jobs�NhK �verbose�K �
warm_start��hN�max_samples�NhhhNhKhKhG        h�auto�hNhG        hG        �feature_names_in_��numpy.core.multiarray��_reconstruct����numpy��ndarray���K ��Cb���R�(KK��h)�dtype����O8�����R�(K�|�NNNJ����J����K?t�b�]�(�Pclass��Sex��Age��SibSp��Parch��Fare��Embarked�et�b�n_features_in_�K�
n_outputs_�K�classes_�h(h+K ��h-��R�(KK��h2�i8�����R�(K�<�NNNJ����J����K t�b�C               �t�b�
n_classes_�K�base_estimator_�h	�estimators_�]�(h)��}�(hhhhhNhKhKhG        hh$hNhJ�
hG        hNhG        hAKhBKhCh(h+K ��h-��R�(KK��h2�f8�����R�(KhKNNNJ����J����K t�b�C              �?�t�bhOh&�scalar���hJC       ���R��max_features_�K�tree_��sklearn.tree._tree��Tree���Kh(h+K ��h-��R�(KK��hJ�C       �t�bK��R�}�(hK�
node_count�M�nodes�h(h+K ��h-��R�(KM��h2�V56�����R�(Kh6N(�
left_child��right_child��feature��	threshold��impurity��n_node_samples��weighted_n_node_samples�t�}�(h{hJK ��h|hJK��h}hJK��h~h[K��hh[K ��h�hJK(��h�h[K0��uK8KKt�b�Bx=         ~                     @�U�Ň�?�           @�@       ]                    �?�b��@��?�            t@       .                     �?.^�����?�             n@                           �?�gtq���?P            �`@       
                  �>@�<ݚ�?             �O@       	                  Y>@�����H�?             "@                        0C�<@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @                           �?�����H�?             K@                           �?@�0�!��?             A@������������������������       �                     6@                          �O@      �?             (@                          �B@      �?              @������������������������       �                     @������������������������       �                      @������������������������       �                     @������������������������       �        
             4@       -                 03�T@X�<ݚ�?0             R@                           �?������?*            �O@������������������������       �                     0@                          �<@(���@��?            �G@                           7@�q�q�?             @������������������������       �                      @������������������������       �                     @       ,                  i?@���� �?            �D@                        ��$:@�G�z��?             4@������������������������       �                     @                        03k:@     ��?             0@������������������������       �                     @        !                 �|Y=@�n_Y�K�?	             *@������������������������       �                     �?"       )                   �J@�q�q�?             (@#       (                   �=@�<ݚ�?             "@$       '                 `f�;@�q�q�?             @%       &                 X��B@z�G�z�?             @������������������������       �      �?              @������������������������       �                     @������������������������       �                     �?������������������������       �                     @*       +                    R@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     5@������������������������       �                     "@/       0                    @Fmq��?F            �Z@������������������������       �                     @1       2                    .@&�����?C            @Y@������������������������       �                     @3       \                    �?L�uϪ�?B            �X@4       E                    �?�Pf����?@            �W@5       6                    �?l��\��?             A@������������������������       �                     @7       D                   �7@ܷ��?��?             =@8       C                    �?�LQ�1	�?             7@9       :                   �9@�C��2(�?             6@������������������������       �      �?              @;       <                   �'@P���Q�?             4@������������������������       �                     @=       >                   �B@      �?
             0@������������������������       �                     $@?       B                   �*@r�q��?             @@       A                    D@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     @������������������������       �                     �?������������������������       �                     @F       [                    �?(��+�?)            �N@G       L                    �?�J�4�?!             I@H       K                 X�l@@      �?             @I       J                 `��,@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @M       N                    >@*
;&���?             G@������������������������       �                     2@O       P                   �?@      �?             <@������������������������       �                     @Q       Z                   @F@���}<S�?             7@R       S                 `fF)@r�q��?
             (@������������������������       �                     @T       Y                   �3@      �?              @U       X                   @D@�q�q�?             @V       W                   �A@z�G�z�?             @������������������������       �      �?              @������������������������       �                     @������������������������       �                     �?������������������������       �                      @������������������������       �                     &@������������������������       �                     &@������������������������       �                     @^       e                    �?H�z���?5             T@_       `                    �?և���X�?             ,@������������������������       �                     @a       b                    �?      �?              @������������������������       �                     @c       d                    5@      �?             @������������������������       �                      @������������������������       �                      @f       u                   �S@�GN�z�?*            �P@g       h                    �?v�X��?             F@������������������������       �                     4@i       j                    �?r�q��?             8@������������������������       �                     @k       n                     �?D�n�3�?             3@l       m                  x�N@z�G�z�?             @������������������������       �                     �?������������������������       �                     @o       t                    �?����X�?	             ,@p       s                    �?�θ�?             *@q       r                   �3@r�q��?             (@������������������������       �                     $@������������������������       �                      @������������������������       �                     �?������������������������       �                     �?v       w                 ���`@�C��2(�?             6@������������������������       �                     "@x       {                 03c@8�Z$���?             *@y       z                 ��)@      �?             @������������������������       �                     @������������������������       �                     �?|       }                   �N@�����H�?             "@������������������������       �                      @������������������������       �                     �?       �                    �?|І"���?�            px@�       �                    �?༉p���?E            �Z@�       �                 pF @>��C��?            �E@�       �                 �|>@ףp=
�?             4@�       �                    �?�}�+r��?             3@������������������������       �                     �?�       �                 �&�@�X�<ݺ?             2@������������������������       �                     �?������������������������       �                     1@������������������������       �                     �?�       �                 ��.@�LQ�1	�?             7@�       �                    �?�<ݚ�?             "@�       �                    @      �?              @������������������������       �                     �?�       �                   �-@؇���X�?             @������������������������       �                     @�       �                 �|Y6@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     �?�       �                 X�,A@@4և���?             ,@������������������������       �                     *@������������������������       �                     �?�       �                 ���1@     ��?(             P@�       �                    @4���C�?            �@@�       �                   �3@     ��?             @@�       �                  �M$@r�q��?             (@������������������������       �                     @�       �                    @���Q��?             @�       �                   �&@      �?             @������������������������       �                      @������������������������       �                      @������������������������       �                     �?�       �                 ���.@���Q��?             4@�       �                   �;@      �?             0@�       �                 pf� @      �?              @�       �                    �?���Q��?             @������������������������       �                     @������������������������       �                      @������������������������       �                     @�       �                    �?      �?              @�       �                 �?� @؇���X�?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @������������������������       �                     �?�       �                   �>@��a�n`�?             ?@�       �                    @ ��WV�?             :@�       �                    @      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     8@�       �                    �?���Q��?             @������������������������       �                      @�       �                   @C@�q�q�?             @������������������������       �                      @������������������������       �                     �?�                          �?�w��.F�?�            �q@�       �                 �?�@�����D�?�            @p@�       �                   �7@     �?Q             `@������������������������       �                     ;@�       �                   �9@���79��??            @Y@�       �                 ���@���Q��?             $@������������������������       �                     @������������������������       �                     @�       �                    �?$�q-�?9            �V@�       �                  s�@$G$n��?            �B@������������������������       �                     0@�       �                 �|Y=@���N8�?             5@������������������������       �                     @�       �                    �?�����H�?
             2@������������������������       �                     @�       �                 �|Y>@"pc�
�?             &@�       �                 ��(@����X�?             @������������������������       ����Q��?             @������������������������       �                      @������������������������       �                     @�       �                   @@@ 7���B�?!             K@�       �                   �?@@-�_ .�?            �B@�       �                 �|Y=@������?             B@������������������������       �                     ,@�       �                  sW@���7�?             6@�       �                 �|�=@�����H�?             "@�       �                 ��,@؇���X�?             @������������������������       �                     @������������������������       �                     �?������������������������       �                      @������������������������       �                     *@������������������������       �                     �?������������������������       �        
             1@�       �                    ,@�`de��?R            �`@������������������������       �                     @�                          �?�+e�X�?M            @_@�       �                    �?0B��D�?H            �]@�       �                    �?      �?             @������������������������       �                     @������������������������       �                     @�       �                 @3�@��Xk�?E             \@�       �                    �?     ��?             0@�       �                    :@�n_Y�K�?             *@������������������������       �                     @�       �                   �A@�����H�?             "@�       �                   �?@      �?             @������������������������       �                     �?������������������������       ��q�q�?             @������������������������       �                     @������������������������       �                     @�                          �?r�q��?=             X@�                          �?p`q�q��?1            �S@�                       `�X#@���y4F�?0             S@�       �                   �3@���}D�?)            �P@�       �                 pf� @�q�q�?             "@�       �                    1@؇���X�?             @������������������������       ��q�q�?             @������������������������       �                     @������������������������       �                      @�       �                   �9@д>��C�?#             M@������������������������       �                     *@�       �                 ��) @�<ݚ�?            �F@�       �                   @F@ȵHPS!�?             :@�       �                   @?@�nkK�?             7@������������������������       �        	             1@�       �                   �@@r�q��?             @������������������������       �                     �?������������������������       �                     @�       �                   �G@�q�q�?             @������������������������       �                      @������������������������       �                     �?                       pf� @p�ݯ��?             3@������������������������       �                     �?                        �?@�q�q�?
             2@                        �;@�eP*L��?             &@������������������������       �                      @                      ���"@X�<ݚ�?             "@������������������������       �                     �?                        �<@      �?              @������������������������       �                      @	      
                �|Y=@�q�q�?             @������������������������       �                     @                      �|�=@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @������������������������       �                     "@������������������������       �                     @������������������������       �                     1@������������������������       �                     @                         �? �q�q�?             8@������������������������       �                     *@                         @�C��2(�?             &@                         @�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                      @�t�b�values�h(h+K ��h-��R�(KMKK��h[�B�        z@     `r@     ``@     �g@     �[@     ``@      G@     @V@      ,@     �H@       @      �?       @      �?       @                      �?      @              @      H@      @      <@              6@      @      @       @      @              @       @              @                      4@      @@      D@      @@      ?@              0@      @@      .@       @      @       @                      @      >@      &@      "@      &@      @              @      &@              @      @       @      �?              @       @       @      @       @      @      �?      @      �?      �?              @      �?                      @       @      �?       @                      �?      5@                      "@      P@      E@      @             �M@      E@              @     �M@     �C@      L@     �C@      @      ?@              @      @      :@      @      4@       @      4@      �?      �?      �?      3@              @      �?      .@              $@      �?      @      �?       @      �?                       @              @      �?                      @     �J@       @      E@       @      @      �?      �?      �?              �?      �?               @             �C@      @      2@              5@      @              @      5@       @      $@       @      @              @       @      @       @      @      �?      �?      �?      @                      �?       @              &@              &@              @              5@     �M@      @       @              @      @       @      @               @       @               @       @              .@     �I@      *@      ?@              4@      *@      &@      @               @      &@      @      �?              �?      @              @      $@      @      $@       @      $@              $@       @              �?              �?               @      4@              "@       @      &@      �?      @              @      �?              �?       @               @      �?             �q@      Z@      J@     �K@      $@     �@@       @      2@      �?      2@              �?      �?      1@      �?                      1@      �?               @      .@      @       @      @       @              �?      @      �?      @              �?      �?              �?      �?              �?              �?      *@              *@      �?              E@      6@      ,@      3@      ,@      2@       @      $@              @       @      @       @       @       @                       @              �?      (@       @      (@      @      @      @       @      @              @       @              @              @      �?      @      �?      @                      �?      �?                      @              �?      <@      @      9@      �?      �?      �?      �?                      �?      8@              @       @       @              �?       @               @      �?             `m@     �H@     �j@      H@     @]@      &@      ;@             �V@      &@      @      @              @      @              U@      @      @@      @      0@              0@      @              @      0@       @      @              "@       @      @       @      @       @       @              @              J@       @     �A@       @     �A@      �?      ,@              5@      �?       @      �?      @      �?      @                      �?       @              *@                      �?      1@             �W@     �B@              @     �W@      >@      V@      >@      @      @      @                      @     @U@      ;@      @      &@      @       @      @              �?       @      �?      @              �?      �?       @              @              @      T@      0@     �O@      0@      N@      0@     �I@      0@      @      @      �?      @      �?       @              @       @              H@      $@      *@             �A@      $@      7@      @      6@      �?      1@              @      �?              �?      @              �?       @               @      �?              (@      @              �?      (@      @      @      @               @      @      @      �?              @      @       @               @      @              @       @      �?       @                      �?      @              "@              @              1@              @              7@      �?      *@              $@      �?       @      �?              �?       @               @        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh$hNhJ/��hG        hNhG        hAKhBKhCh(h+K ��h-��R�(KK��h[�C              �?�t�bhOh`hJC       ���R�hdKhehhKh(h+K ��h-��R�(KK��hJ�C       �t�bK��R�}�(hKhrM#hsh(h+K ��h-��R�(KM#��hz�B�?         &                   �1@�)�>_M�?�           @�@                           @��>4և�?4             U@       
                     @���!pc�?(            �P@                           �?�C��2(�?            �@@������������������������       �        	             0@                        ���`@@�0�!��?
             1@������������������������       �                     (@       	                 �(\�?���Q��?             @������������������������       �                      @������������������������       �                     @                          �,@�eP*L��?            �@@                        `��+@�r����?
             .@������������������������       �                     @                          �3@      �?              @                          �/@�q�q�?             @������������������������       �                     �?                           @      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @                        pf� @�E��ӭ�?             2@                           �?      �?             $@                           �?r�q��?             @������������������������       �                     @������������������������       �      �?              @������������������������       �                     @������������������������       �                      @                           @r�q��?             2@������������������������       �                     @                           �?d}h���?	             ,@������������������������       �                     @        %                 ���A@���!pc�?             &@!       "                 ��T?@և���X�?             @������������������������       �                      @#       $                    @���Q��?             @������������������������       �                     @������������������������       �                      @������������������������       �                     @'       ~                    �?J�
��O�?�           ��@(       ?                     @���*�?y            @h@)       0                    �?Hn�.P��?H             _@*       /                   �*@��v$���?&            �N@+       ,                   �'@�X�<ݺ?             2@������������������������       �                     @-       .                    ;@�C��2(�?             &@������������������������       �      �?              @������������������������       �                     "@������������������������       �                    �E@1       <                    �?�[|x��?"            �O@2       ;                    �?      �?             H@3       4                   �6@=QcG��?            �G@������������������������       �                      @5       :                    :@����?�?            �F@6       7                    �?�C��2(�?             &@������������������������       �                      @8       9                    D@�����H�?             "@������������������������       �                      @������������������������       �                     �?������������������������       �                     A@������������������������       �                     �?=       >                 ���`@�r����?             .@������������������������       �                     *@������������������������       �                      @@       i                    �?��(@��?1            �Q@A       L                    �?\X��t�?!             G@B       I                 pF @�z�G��?             4@C       F                 ���@؇���X�?
             ,@D       E                    �?�q�q�?             @������������������������       �                      @������������������������       �                     �?G       H                 �|>@�C��2(�?             &@������������������������       �                     $@������������������������       �                     �?J       K                 ���2@�q�q�?             @������������������������       �                     @������������������������       �                      @M       T                   �@��
ц��?             :@N       Q                 pff@      �?              @O       P                 �|�9@      �?              @������������������������       �                     �?������������������������       �                     �?R       S                   �<@r�q��?             @������������������������       �                     @������������������������       �                     �?U       h                    �?�q�q�?             2@V       Y                    3@ҳ�wY;�?             1@W       X                 `F�+@�q�q�?             @������������������������       �                      @������������������������       �                     �?Z       a                    �?����X�?	             ,@[       `                 pf� @�����H�?             "@\       ]                 �?�@z�G�z�?             @������������������������       �                     @^       _                    9@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @b       c                 �|Y>@���Q��?             @������������������������       �                      @d       e                   �@@�q�q�?             @������������������������       �                     �?f       g                   �D@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     �?j       w                 �A7@�q�q�?             8@k       r                    �?      �?	             $@l       m                    5@      �?             @������������������������       �                     �?n       q                   �/@���Q��?             @o       p                    �?�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                      @s       t                    �?      �?             @������������������������       �                     �?u       v                 032@�q�q�?             @������������������������       �                      @������������������������       �                     �?x       y                 ��A>@؇���X�?             ,@������������������������       �                     @z       }                    �?����X�?             @{       |                    @�q�q�?             @������������������������       �                     @������������������������       �                      @������������������������       �                     �?       �                     �?�*�@P��?            {@�       �                    �?�lg����?7            �U@�       �                    �?L
�q��?(            �M@�       �                 �|�;@������?             1@������������������������       �                      @�       �                 p�w@�r����?             .@�       �                   �J@@4և���?             ,@������������������������       �                      @�       �                   �L@r�q��?             @�       �                  ��@@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @������������������������       �                     �?�       �                   @@@�ՙ/�?             E@�       �                    �?r�q��?             2@�       �                 `fF<@@�0�!��?
             1@�       �                 `fF:@և���X�?             @������������������������       �                     @�       �                 �|�<@      �?             @������������������������       �                      @������������������������       �      �?              @������������������������       �                     $@������������������������       �                     �?�       �                   �J@r�q��?             8@�       �                   �9@8�Z$���?             *@������������������������       �                     �?�       �                    G@�8��8��?             (@������������������������       �                     @�       �                   �D@z�G�z�?             @������������������������       �                     @������������������������       �                     �?�       �                 `fF<@"pc�
�?             &@������������������������       �                     @�       �                   @>@�q�q�?             @������������������������       �                      @������������������������       �                     @�       �                    �?X�<ݚ�?             ;@�       �                 ��sW@r�q��?             @������������������������       �                     @������������������������       �                     �?�       �                    �?�q�q�?             5@������������������������       �                     @�       �                    �?b�2�tk�?
             2@�       �                    �?��S���?	             .@�       �                  x#J@և���X�?             ,@������������������������       �                     @�       �                 `�iJ@���Q��?             $@������������������������       �                     @�       �                 03�S@և���X�?             @�       �                    <@z�G�z�?             @������������������������       �                     �?������������������������       �                     @������������������������       �                      @������������������������       �                     �?������������������������       �                     @�       �                     @�:���?�            �u@�       �                    9@��?^�k�?-            �Q@������������������������       �        #            �J@�       �                    @@�t����?
             1@�       �                   �H@      �?              @������������������������       �                      @������������������������       �                     @������������������������       �                     "@�       �                 �?�@��l�5�?�            `q@�       �                    �?,_ʯ08�?`            �c@�       �                 �{@��4@��?^            @c@�       �                    �?�X�C�?E             \@�       �                  ��@ �h�7W�?!            �J@�       �                   �7@������?             B@�       �                   �5@r�q��?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     >@�       �                 �|Y>@�t����?             1@������������������������       �r�q��?             (@������������������������       �                     @�       �                 �?$@�:�B��?$            �M@�       �                 �|�=@���H��?             E@�       �                    7@z�G�z�?             9@������������������������       �                     "@�       �                   �9@     ��?             0@�       �                 `fF@      �?              @�       �                   �8@z�G�z�?             @�       �                 �&b@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                      @������������������������       �                     @�       �                 ��,@      �?              @������������������������       �                     @�       �                 �|�;@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     1@�       �                    >@�t����?	             1@�       �                   �9@z�G�z�?             .@������������������������       �                     @�       �                   �;@      �?              @������������������������       �                     @������������������������       �                     @������������������������       �                      @������������������������       �                     E@������������������������       �                     @�       �                   �4@�O��=�?M            �]@�       �                    �?��S���?
             .@�       �                   �3@���|���?             &@�       �                 ��Y @և���X�?             @������������������������       �                     @������������������������       �                     @������������������������       �                     @�       �                    �?      �?             @������������������������       �                      @�       �                 8#�1@      �?              @������������������������       �                     �?������������������������       �                     �?�                          @F@D>�Q�?C             Z@�                         @@@�+�ԗ�??            �X@�                          �?$]��<C�?/            �Q@�                       ��q1@�*/�8V�?            �G@�       �                    �?� ��1�?            �D@������������������������       �                     �?�                         �>@z�G�z�?             D@�       �                 ��) @��� ��?             ?@������������������������       �        
             3@�       �                 ��� @�q�q�?	             (@������������������������       �                      @�                         @=@z�G�z�?             $@�                          �8@�����H�?             "@������������������������       �                     @                      ��)"@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     �?                      @3�@X�<ݚ�?             "@                        �?@�q�q�?             @������������������������       �                     �?������������������������       �z�G�z�?             @	      
                ��i @�q�q�?             @������������������������       �                      @������������������������       �                     �?                         ;@�q�q�?             @������������������������       �                     �?                      �|�<@���Q��?             @������������������������       �                     �?                      �|�>@      �?             @������������������������       ��q�q�?             @������������������������       �                     �?                      ��.@�8��8��?             8@                         �?����X�?             @                      �|Y<@�q�q�?             @������������������������       �                     @������������������������       �                      @������������������������       �                     �?������������������������       �                     1@                        �E@ 7���B�?             ;@������������������������       �                     5@                         �?r�q��?             @                      @3�@      �?             @������������������������       �                     �?������������������������       �                     @������������������������       �                      @!      "                   G@      �?             @������������������������       �                     @������������������������       �                     @�t�bh�h(h+K ��h-��R�(KM#KK��h[�B0       `{@      q@     �@@     �I@      2@      H@      @      >@              0@      @      ,@              (@      @       @               @      @              .@      2@       @      *@              @       @      @       @      �?      �?              �?      �?              �?      �?                      @      *@      @      @      @      �?      @              @      �?      �?      @               @              .@      @      @              &@      @      @               @      @      @      @       @               @      @              @       @              @             Py@     �k@     �E@     �b@      @     �]@      �?      N@      �?      1@              @      �?      $@      �?      �?              "@             �E@      @      M@      @     �F@      @      F@       @              �?      F@      �?      $@               @      �?       @               @      �?                      A@              �?       @      *@              *@       @             �B@     �@@      4@      :@      @      ,@       @      (@      �?       @               @      �?              �?      $@              $@      �?              @       @      @                       @      ,@      (@       @      @      �?      �?              �?      �?              �?      @              @      �?              (@      @      &@      @      �?       @               @      �?              $@      @       @      �?      @      �?      @              �?      �?      �?                      �?      @               @      @               @       @      �?      �?              �?      �?              �?      �?              �?              1@      @      @      @      @      @      �?               @      @       @      �?       @                      �?               @       @       @              �?       @      �?       @                      �?      (@       @      @              @       @      @       @      @                       @      �?             �v@      R@      K@      @@     �C@      4@      *@      @               @      *@       @      *@      �?       @              @      �?      �?      �?      �?                      �?      @                      �?      :@      0@      .@      @      ,@      @      @      @      @              �?      @               @      �?      �?      $@              �?              &@      *@       @      &@      �?              �?      &@              @      �?      @              @      �?              "@       @      @              @       @               @      @              .@      (@      �?      @              @      �?              ,@      @      @              &@      @       @      @       @      @      @              @      @              @      @      @      @      �?              �?      @                       @              �?      @             @s@      D@      Q@       @     �J@              .@       @      @       @               @      @              "@              n@      C@     @b@      *@     �a@      *@     �X@      *@      I@      @     �A@      �?      @      �?      @                      �?      >@              .@       @      $@       @      @             �H@      $@     �B@      @      4@      @      "@              &@      @      @      @      �?      @      �?       @      �?                       @               @      @              @      �?      @               @      �?       @                      �?      1@              (@      @      (@      @      @              @      @              @      @                       @      E@              @             �W@      9@       @      @      @      @      @      @              @      @              @              �?      @               @      �?      �?              �?      �?             �U@      2@     �T@      .@     �L@      ,@     �A@      (@     �@@       @      �?              @@       @      ;@      @      3@               @      @               @       @       @       @      �?      @               @      �?              �?       @                      �?      @      @      @       @              �?      @      �?      �?       @               @      �?               @      @              �?       @      @      �?              �?      @      �?       @              �?      6@       @      @       @      @       @      @                       @      �?              1@              :@      �?      5@              @      �?      @      �?              �?      @               @              @      @              @      @        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh$hNhJu�7hG        hNhG        hAKhBKhCh(h+K ��h-��R�(KK��h[�C              �?�t�bhOh`hJC       ���R�hdKhehhKh(h+K ��h-��R�(KK��hJ�C       �t�bK��R�}�(hKhrM)hsh(h+K ��h-��R�(KM)��hz�B�@         "                   @^80�B�?�           @�@       �                    �?��E�Ϩ�?�           `�@       8                    �?�H&��?<           `~@                            @nS�2ִ�?]            �`@                          �*@��pBI�?1            @R@                          �B@�KM�]�?             3@       
                   �9@��S�ۿ?
             .@       	                   �6@؇���X�?             @������������������������       �                     @������������������������       �      �?              @������������������������       �                      @                          �'@      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �        %             K@                           �?�p����?,            �N@                           0@և���X�?             @������������������������       �                      @                           �?z�G�z�?             @������������������������       �                     @                         S�2@      �?              @������������������������       �                     �?������������������������       �                     �?       )                 �̌@���3L�?&             K@                            �?�z�G��?             >@                        �|>@�d�����?             3@                           �?      �?             0@                        ���@��S�ۿ?             .@������������������������       �                     �?������������������������       �                     ,@������������������������       �                     �?������������������������       �                     @!       "                 ���@���|���?             &@������������������������       �                     @#       &                 �&B@�q�q�?             @$       %                   �7@      �?             @������������������������       �                     �?������������������������       �                     @'       (                   �<@      �?              @������������������������       �                     �?������������������������       �                     �?*       7                   �;@�q�q�?             8@+       6                   �7@      �?             0@,       5                    3@�eP*L��?             &@-       .                    �?����X�?             @������������������������       �                      @/       4                    ,@���Q��?             @0       1                    �?�q�q�?             @������������������������       �                     �?2       3                    @      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @������������������������       �                     @������������������������       �                     @������������������������       �                      @9       �                 ��$:@�g���E�?�             v@:       ;                    $@�S</�z�?�            `q@������������������������       �                     @<       g                 �|Y=@�u����?�             q@=       F                    �?�>4և��?F             \@>       ?                     @�q�q�?             (@������������������������       �                     �?@       A                 �Y�@�eP*L��?             &@������������������������       �                     @B       E                    �?����X�?             @C       D                   �2@      �?             @������������������������       �                      @������������������������       �                      @������������������������       �                     @G       ^                 ��Y @R���Q�?@             Y@H       Y                 @3�@Z���c��?)            �O@I       L                 ���@8�Z$���?              J@J       K                 ���@�q�q�?             (@������������������������       �                      @������������������������       �                     @M       N                 �?$@ףp=
�?             D@������������������������       �        
             .@O       X                 �1@�J�4�?             9@P       Q                   �3@���Q��?             $@������������������������       �                     @R       W                   �;@�q�q�?             @S       T                   �6@z�G�z�?             @������������������������       �                      @U       V                   �9@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     �?������������������������       �                     .@Z       ]                   �3@�eP*L��?	             &@[       \                    1@r�q��?             @������������������������       ��q�q�?             @������������������������       �                     @������������������������       �                     @_       f                   �3@@-�_ .�?            �B@`       a                   �2@؇���X�?
             ,@������������������������       �                     $@b       e                     @      �?             @c       d                   �'@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     �?������������������������       �                     7@h       �                    �?xdQ�m��?h            @d@i       �                   @@@���`uӽ?g             d@j       {                   �?@<����?<            �W@k       v                 ��) @���1j	�?5            �U@l       m                  s�@��.N"Ҭ?,            @Q@������������������������       �                    �@@n       o                    �?�X�<ݺ?             B@������������������������       �                     @p       u                 �|�=@�FVQ&�?            �@@q       r                    �?�>����?             ;@������������������������       �ףp=
�?             $@s       t                  sW@�IєX�?
             1@������������������������       �      �?             @������������������������       �                     *@������������������������       �                     @w       x                    �?@�0�!��?	             1@������������������������       �                      @y       z                 �̜"@��S�ۿ?             .@������������������������       �                     �?������������������������       �                     ,@|       }                     @�q�q�?             "@������������������������       �                     �?~                        P�@      �?              @������������������������       �                     �?�       �                 @3�@����X�?             @������������������������       �z�G�z�?             @�       �                 ��i @      �?              @������������������������       �                     �?������������������������       �                     �?�       �                 �?�@Pa�	�?+            �P@������������������������       �                     <@�       �                     @�}�+r��?             C@�       �                   @F@XB���?             =@�       �                   @D@��S�ۿ?	             .@������������������������       �                     *@������������������������       �      �?              @������������������������       �                     ,@�       �                 @3�@�����H�?             "@�       �                   �D@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @������������������������       �                     �?�       �                    �?` .�(�?/            �R@�       �                 ��";@���Q��?+            �Q@�       �                 03k:@8����?
             7@������������������������       �                     @�       �                   @L@b�2�tk�?             2@�       �                   @G@������?             .@�       �                 X��B@���|���?             &@�       �                 �|�<@      �?              @������������������������       �                     @������������������������       �z�G�z�?             @������������������������       �                     @������������������������       �                     @������������������������       �                     @�       �                    �?�*/�8V�?!            �G@�       �                    �?�(�Tw��?            �C@�       �                 p�i@@�q�q�?	             (@�       �                   �<@      �?              @������������������������       �                     @������������������������       �                     @������������������������       �                     @�       �                 0�K@�<ݚ�?             ;@�       �                   @>@ףp=
�?             4@�       �                   `O@����X�?             @������������������������       �                     @������������������������       �                      @������������������������       �        
             *@�       �                   �7@և���X�?             @������������������������       �                     �?�       �                 lfda@�q�q�?             @�       �                 �|�;@z�G�z�?             @������������������������       �                     @�       �                 �|�>@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     �?�       �                    �?      �?              @�       �                   @B@z�G�z�?             @�       �                    >@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @������������������������       �                     @�       �                    ?@      �?             @������������������������       �                     @������������������������       �                     �?�                          @�'�=z��?            �h@�       �                     @rѱ�D��?w            �f@�       �                    �?tp�P�?G            @[@�       �                 �|�=@��}*_��?             ;@������������������������       �        	             &@�       �                   �A@      �?
             0@������������������������       �                     @�       �                    �?���Q��?             $@������������������������       �                     @�       �                    �?z�G�z�?             @�       �                 �UkT@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @�       �                    �?�4F����?4            �T@�       �                    �?�:�^���?            �F@�       �                    E@�X�<ݺ?             B@�       �                     �?XB���?             =@������������������������       �                     (@�       �                    �?�IєX�?
             1@�       �                    �?      �?	             0@�       �                   �7@ףp=
�?             $@������������������������       �                     �?������������������������       �                     "@������������������������       �                     @������������������������       �                     �?�       �                     �?؇���X�?             @������������������������       �                     @������������������������       �                     �?�       �                 ���`@�<ݚ�?             "@������������������������       �                     @������������������������       �                      @�       �                    -@�Gi����?            �B@������������������������       �                     "@�       �                     �?d}h���?             <@�       �                    �?և���X�?
             ,@�       �                    G@�n_Y�K�?	             *@�       �                    �?      �?             $@�       �                  x#J@X�<ݚ�?             "@������������������������       �                      @�       �                    >@և���X�?             @������������������������       �                      @�       �                 `f�K@z�G�z�?             @�       �                   �C@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @������������������������       �                     �?������������������������       �                     @������������������������       �                     �?������������������������       �                     ,@�       �                  S�$@X~�pX��?0            @R@�       �                    �?�C��2(�?             &@������������������������       �                     �?�       �                 �&B@ףp=
�?             $@������������������������       �                     @�       �                    4@z�G�z�?             @������������������������       �                     �?������������������������       �                     @�       �                 ��Y)@f���M�?(             O@������������������������       �                     @�                          �?��U/��?%            �L@�                       `v�6@`��}3��?!            �J@�                          /@Z�K�D��?            �G@                          �?���!pc�?             &@                       S%/@�z�G��?             $@                      03�-@և���X�?             @                        �-@�q�q�?             @������������������������       �                      @������������������������       �                     @������������������������       �                     �?������������������������       �                     @������������������������       �                     �?	                      �q5@      �?             B@
                      �?�-@H�V�e��?             A@������������������������       �                     &@                         �?8����?             7@                      ���/@����X�?             @                         �?�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     @                      �|�<@      �?             0@������������������������       �                     @                      �|�>@r�q��?
             (@                         �?      �?              @������������������������       �                     @������������������������       �                      @������������������������       �                     @������������������������       �                      @������������������������       �                     @������������������������       �                     @                        @C@      �?             0@                         �?z�G�z�?             @������������������������       �                     @������������������������       �                     �?       !                    @"pc�
�?             &@������������������������       �                      @������������������������       �                     "@#      (                   �?h�����?             <@$      %                   �?$�q-�?	             *@������������������������       �                     @&      '                ���d@�����H�?             "@������������������������       �                      @������������������������       �                     �?������������������������       �                     .@�t�bh�h(h+K ��h-��R�(KM)KK��h[�B�       p{@     q@     �y@      q@     �s@     @e@      =@     @Z@       @     �Q@       @      1@      �?      ,@      �?      @              @      �?      �?               @      �?      @              @      �?                      K@      ;@      A@      @      @               @      @      �?      @              �?      �?      �?                      �?      7@      ?@      "@      5@      @      ,@       @      ,@      �?      ,@      �?                      ,@      �?              @              @      @              @      @       @      @      �?              �?      @              �?      �?              �?      �?              ,@      $@      @      $@      @      @       @      @               @       @      @       @      �?      �?              �?      �?              �?      �?                       @      @                      @       @             �q@     @P@     �n@      A@              @     �n@      >@      W@      4@      @      @      �?              @      @      @               @      @       @       @       @                       @              @     @U@      .@      I@      *@      F@       @       @      @       @                      @      B@      @      .@              5@      @      @      @      @               @      @      �?      @               @      �?       @      �?                       @      �?              .@              @      @      �?      @      �?       @              @      @             �A@       @      (@       @      $@               @       @      �?       @               @      �?              �?              7@              c@      $@     �b@      $@     �U@       @     @T@      @     �P@       @     �@@              A@       @      @              ?@       @      9@       @      "@      �?      0@      �?      @      �?      *@              @              ,@      @               @      ,@      �?              �?      ,@              @      @      �?              @      @              �?      @       @      @      �?      �?      �?              �?      �?              P@       @      <@              B@       @      <@      �?      ,@      �?      *@              �?      �?      ,@               @      �?      �?      �?      �?                      �?      @              �?             �E@      ?@      E@      <@      @      0@              @      @      &@      @      &@      @      @      �?      @              @      �?      @      @                      @      @             �A@      (@      <@      &@      @      @      @      @      @                      @      @              5@      @      2@       @      @       @      @                       @      *@              @      @      �?               @      @      �?      @              @      �?      �?      �?                      �?      �?              @      �?      @      �?      �?      �?      �?                      �?      @              @              �?      @              @      �?              X@     �Y@     �U@      X@      B@     @R@      $@      1@              &@      $@      @      @              @      @              @      @      �?      �?      �?              �?      �?              @              :@      L@      @     �D@       @      A@      �?      <@              (@      �?      0@      �?      .@      �?      "@      �?                      "@              @              �?      �?      @              @      �?               @      @              @       @              6@      .@              "@      6@      @       @      @       @      @      @      @      @      @       @              @      @       @              �?      @      �?      �?      �?                      �?              @              �?      @                      �?      ,@              I@      7@      $@      �?      �?              "@      �?      @              @      �?              �?      @              D@      6@              @      D@      1@      B@      1@      >@      1@      @       @      @      @      @      @       @      @       @                      @      �?                      @              �?      ;@      "@      ;@      @      &@              0@      @       @      @       @      �?              �?       @                      @      ,@       @      @              $@       @      @       @      @                       @      @                       @      @              @              $@      @      �?      @              @      �?              "@       @               @      "@              ;@      �?      (@      �?      @               @      �?       @                      �?      .@        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh$hNhJ��!XhG        hNhG        hAKhBKhCh(h+K ��h-��R�(KK��h[�C              �?�t�bhOh`hJC       ���R�hdKhehhKh(h+K ��h-��R�(KK��hJ�C       �t�bK��R�}�(hKhrMEhsh(h+K ��h-��R�(KME��hz�BG         �                 �J/@^IB�A��?�           @�@                           /@���!pc�?�            x@                        P��%@ףp=
�?             4@                           �?����X�?             @������������������������       �                     @������������������������       �                      @������������������������       �                     *@       �                   @@@�8��<�?�            �v@	       0                    �?,�?���?�            �q@
                          �0@�����?4            �S@������������������������       �                      @                           �?*-ڋ�p�?2            @S@                           �?�+$�jP�?             ;@                           4@���Q��?             @������������������������       �                     �?                           �?      �?             @                        ��	-@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @                           �?��2(&�?             6@                        pF @P���Q�?             4@������������������������       �        
             .@                           �?z�G�z�?             @                            @      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @       %                  ��@�J�4�?             I@       $                   �6@��S�ۿ?             >@        #                    �?����X�?             @!       "                    5@���Q��?             @������������������������       �                     @������������������������       �                      @������������������������       �                      @������������������������       �                     7@&       )                    �?�z�G��?             4@'       (                    �?      �?             @������������������������       �                     @������������������������       �                     @*       /                   @'@d}h���?
             ,@+       ,                 �|Y=@�z�G��?             $@������������������������       �                      @-       .                 �|Y>@      �?              @������������������������       �r�q��?             @������������������������       �                      @������������������������       �                     @1       |                 �|Y=@�Ј� �?�            �i@2       i                   �:@4kMU*m�?X            `a@3       h                    �?,y�xEE�?D            �Z@4       a                   �8@ ��/K��?C            �Z@5       R                 0S5 @jJA��v�?7            �V@6       7                    1@T����1�?#             M@������������������������       ��q�q�?             @8       =                   �2@�2�o�U�?!            �K@9       <                    �?      �?              @:       ;                 ��@؇���X�?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     �?>       I                 �1@"Ae���?            �G@?       @                    �?П[;U��?             =@������������������������       �                      @A       F                 �?$@���N8�?             5@B       C                    7@�t����?
             1@������������������������       �                     ,@D       E                 �&b@�q�q�?             @������������������������       �                     �?������������������������       �                      @G       H                   �6@      �?             @������������������������       �                     @������������������������       �                     �?J       Q                    �?r�q��?             2@K       L                    �?�t����?             1@������������������������       �                     �?M       N                 @3�@      �?             0@������������������������       �                     $@O       P                   �3@�q�q�?             @������������������������       �                      @������������������������       �                     @������������������������       �                     �?S       ^                   �7@�C��2(�?            �@@T       U                 @�"@`Jj��?             ?@������������������������       �                     &@V       W                 ���"@ףp=
�?             4@������������������������       �                     �?X       ]                    �?�}�+r��?             3@Y       Z                   �4@�IєX�?	             1@������������������������       �                     (@[       \                 pF%@z�G�z�?             @������������������������       �                     �?������������������������       �                     @������������������������       �                      @_       `                     @      �?              @������������������������       �                     �?������������������������       �                     �?b       g                    �?��S�ۿ?             .@c       f                    �?�q�q�?             @d       e                 pff@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     �?������������������������       �        	             (@������������������������       �                     �?j       {                    �?     ��?             @@k       l                    �?`՟�G��?             ?@������������������������       �                     "@m       t                   �;@�GN�z�?             6@n       o                     @      �?              @������������������������       �                     @p       q                 pb@���Q��?             @������������������������       �                      @r       s                 �� @�q�q�?             @������������������������       �                      @������������������������       �                     �?u       v                   �<@؇���X�?
             ,@������������������������       �                     @w       x                 ���"@      �?              @������������������������       �                     @y       z                     @      �?             @������������������������       �                      @������������������������       �                      @������������������������       �                     �?}       �                   �>@�� =[�?)             Q@~       �                 �|�=@ףp=
�?              I@       �                    �?�KM�]�?             C@������������������������       �                      @�       �                 ��) @�����H�?             B@�       �                  sW@`Jj��?             ?@�       �                     @8�Z$���?	             *@������������������������       �                     @�       �                 ��,@����X�?             @������������������������       �                     @������������������������       �      �?             @������������������������       �                     2@�       �                     @���Q��?             @������������������������       �                     �?�       �                 �̜!@      �?             @������������������������       �                     �?������������������������       �                     @�       �                     @�8��8��?             (@������������������������       �                     @�       �                 �̌!@�����H�?             "@������������������������       �                      @������������������������       �                     �?�       �                    �?�q�q�?	             2@�       �                 ج�$@�q�q�?             @������������������������       �                     @������������������������       �                      @�       �                   �?@�q�q�?             (@������������������������       �                      @�       �                 P�@z�G�z�?             $@������������������������       �                     �?�       �                     @�����H�?             "@������������������������       �                      @�       �                 @3�@؇���X�?             @������������������������       �                     @�       �                 ��i @      �?              @������������������������       �                     �?������������������������       �                     �?�       �                 �?�@l{��b��?5            �S@������������������������       �                     @@�       �                    �?��E�B��?            �G@�       �                   �'@�q�q�?             @������������������������       �                     @�       �                   �B@�q�q�?             @������������������������       �                     �?������������������������       �                      @�       �                 pFt @������?            �D@�       �                    �?z�G�z�?             $@�       �                   �E@�<ݚ�?             "@������������������������       �                     @�       �                   �G@      �?             @������������������������       �                      @������������������������       �                      @������������������������       �                     �?������������������������       �                     ?@�                            @��e��?�            pt@�                          @$��m��?�            @m@�       
                   �?X������?�             m@�       �                    �?`��2�i�?�            �i@�       �                    �?�c:��?>             W@�       �                    �?���7�?             F@�       �                   �G@�C��2(�?             6@������������������������       �                     1@�       �                 ��-K@���Q��?             @������������������������       �                      @������������������������       �                     @������������������������       �                     6@�       �                     �?8��8���?!             H@������������������������       �                     :@�       �                   �7@�GN�z�?             6@������������������������       �                      @�       �                    �?R���Q�?             4@�       �                  	<@�z�G��?             $@�       �                    D@�q�q�?             "@������������������������       �                     @������������������������       �                     @������������������������       �                     �?������������������������       �                     $@�       �                    �?>4և���?M             \@�       �                 �D@E@��7��?+            �N@�       �                    �?�p ��?            �D@�       �                    �?      �?             D@�       �                 X�,@@���Q��?             $@�       �                 0C�<@z�G�z�?             @������������������������       �                     @������������������������       �                     �?�       �                 `v�<@���Q��?             @������������������������       �                      @�       �                   �O@�q�q�?             @�       �                  ��@@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     �?�       �                   �J@��S���?             >@�       �                 ��$:@�q�q�?             8@������������������������       �                     @�       �                   �E@�S����?             3@�       �                 �|�?@$�q-�?	             *@�       �                 `f�<@r�q��?             @�       �                 �|�<@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @������������������������       �                     @�       �                   �G@�q�q�?             @�       �                  I>@      �?             @������������������������       ��q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     @������������������������       �                     �?�       �                 �̾w@R���Q�?             4@������������������������       �                     1@������������������������       �                     @�       �                    <@��e�B��?"            �I@�       �                 h"P@�t����?             1@�       �                    �?      �?             0@�       �                    6@؇���X�?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     "@������������������������       �                     �?�       �                  x#J@������?             A@�       �                    :@�8��8��?             (@�       �                   �@@z�G�z�?             @�       �                    �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @������������������������       �                     @�       �                 `�iJ@�X����?             6@������������������������       �                      @                          �?      �?             4@                      @�pX@և���X�?             @������������������������       �                     @������������������������       �                     @      	                   �?$�q-�?             *@                        �B@ףp=
�?             $@������������������������       �                     @                        �D@z�G�z�?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     @                         @>���Rp�?             =@                         �?      �?             <@                          �?�r����?             .@                         �?z�G�z�?             $@������������������������       �                     @                          @����X�?             @������������������������       �                     �?                      ���`@r�q��?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     @                          �?�n_Y�K�?	             *@                         6@z�G�z�?             @������������������������       �                     @������������������������       �                     �?                         �?      �?              @                        �;@z�G�z�?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     @������������������������       �                     �?������������������������       �                     �?!      .                @3�4@<)�%�w�?:            @W@"      '                   �?�P�*�?             ?@#      &                �|�7@�����H�?             "@$      %                   �?      �?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     @(      )                   �?�eP*L��?             6@������������������������       �                     @*      -                   �?      �?             0@+      ,                   +@�	j*D�?
             *@������������������������       �                     @������������������������       �                     "@������������������������       �                     @/      8                   �?t�7��?'             O@0      1                �T)D@���Q��?	             .@������������������������       �                     @2      3                   ;@�q�q�?             "@������������������������       �                     �?4      5                �|�<@      �?              @������������������������       �                     �?6      7                �|�>@����X�?             @������������������������       ��q�q�?             @������������������������       �                     �?9      :                   �?�*/�8V�?            �G@������������������������       �                      @;      @                   @��S�ۿ?            �F@<      =                   �?"pc�
�?             &@������������������������       �                     @>      ?                   @      �?             @������������������������       �                      @������������������������       �                      @A      B                   @г�wY;�?             A@������������������������       �                     =@C      D                ��T?@z�G�z�?             @������������������������       �                     @������������������������       �                     �?�t�b��     h�h(h+K ��h-��R�(KMEKK��h[�BP       �z@     �q@     �q@     @Z@       @      2@       @      @              @       @                      *@     `q@     �U@     �i@     @T@     �G@      @@               @     �G@      >@      @      6@       @      @      �?              �?      @      �?      �?              �?      �?                       @      @      3@      �?      3@              .@      �?      @      �?      @              @      �?                      �?       @              E@       @      <@       @      @       @      @       @      @                       @       @              7@              ,@      @      @      @      @                      @      &@      @      @      @               @      @      �?      @      �?       @              @             �c@     �H@     @Y@      C@     �T@      8@     �T@      7@     @Q@      6@     �C@      3@      �?       @      C@      1@      @      �?      @      �?      @                      �?      �?              ?@      0@      0@      *@               @      0@      @      .@       @      ,@              �?       @      �?                       @      �?      @              @      �?              .@      @      .@       @      �?              ,@       @      $@              @       @               @      @                      �?      >@      @      =@       @      &@              2@       @              �?      2@      �?      0@      �?      (@              @      �?              �?      @               @              �?      �?              �?      �?              ,@      �?       @      �?      �?      �?      �?                      �?      �?              (@                      �?      2@      ,@      1@      ,@              "@      1@      @      @      @      @               @      @               @       @      �?       @                      �?      (@       @      @              @       @      @               @       @       @                       @      �?             �L@      &@     �F@      @      A@      @       @              @@      @      =@       @      &@       @      @              @       @      @               @       @      2@              @       @              �?      @      �?              �?      @              &@      �?      @               @      �?       @                      �?      (@      @      @       @      @                       @       @      @               @       @       @              �?       @      �?       @              @      �?      @              �?      �?              �?      �?             @R@      @      @@             �D@      @       @      @              @       @      �?              �?       @             �C@       @       @       @      @       @      @               @       @               @       @              �?              ?@              b@     �f@     @T@      c@      T@      c@     @R@     ``@      @     @U@       @      E@       @      4@              1@       @      @       @                      @              6@      @     �E@              :@      @      1@       @              @      1@      @      @      @      @              @      @                      �?              $@     �P@      G@      C@      7@      5@      4@      4@      4@      @      @      @      �?      @                      �?       @      @               @       @      �?      �?      �?      �?                      �?      �?              ,@      0@       @      0@      @              @      0@      �?      (@      �?      @      �?       @               @      �?                      @              @       @      @       @       @      �?       @      �?                       @      @              �?              1@      @      1@                      @      <@      7@       @      .@      �?      .@      �?      @      �?                      @              "@      �?              :@       @      &@      �?      @      �?      �?      �?      �?                      �?      @              @              .@      @               @      .@      @      @      @              @      @              (@      �?      "@      �?      @              @      �?              �?      @              @              @      6@      @      5@       @      *@       @       @              @       @      @      �?              �?      @              @      �?                      @      @       @      �?      @              @      �?              @      @      �?      @      �?                      @      @                      �?      �?              P@      =@      *@      2@      �?       @      �?      @      �?                      @              @      (@      $@              @      (@      @      "@      @              @      "@              @             �I@      &@      "@      @      @              @      @              �?      @      @      �?               @      @       @      @              �?      E@      @               @      E@      @      "@       @      @               @       @       @                       @     �@@      �?      =@              @      �?      @                      �?�t�bubhhubh)��}�(hhhhhNhKhKhG        hh$hNhJC�NhG        hNhG        hAKhBKhCh(h+K ��h-��R�(KK��h[�C              �?�t�bhOh`hJC       ���R�hdKhehhKh(h+K ��h-��R�(KK��hJ�C       �t�bK��R�}�(hKhrM+hsh(h+K ��h-��R�(KM+��hz�BhA         �                     @4�<����?�           @�@       	                   �1@��~���?�            �u@                        ���`@�X�<ݺ?             B@������������������������       �                     @@                           �?      �?             @                           �?�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     �?
       S                     �?���>4��?�            @s@                           �?��T���?p            �f@                          �H@`׀�:M�?,            �R@������������������������       �        #             M@                          @I@      �?	             0@������������������������       �                     �?������������������������       �                     .@       R                 �̾w@�W;�E��?D            �Z@       '                    �? s�n_Y�?C             Z@       &                 @�pX@      �?             B@       %                    �?��H�}�?             9@                        ��";@���N8�?             5@������������������������       �                     �?       $                    �?z�G�z�?             4@                           C@������?	             1@                         Y>@�����H�?             "@                        �|�;@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     @       #                   �O@      �?              @       "                   �I@      �?             @        !                 �̌K@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @������������������������       �                     @������������������������       �                     @������������������������       �                     @������������������������       �                     &@(       )                 ��$:@�����?/             Q@������������������������       �                      @*       +                   x:@d��0u��?)             N@������������������������       �                      @,       I                   �E@&y�X���?'             M@-       .                    8@�4�����?             ?@������������������������       �                     @/       F                    �?X�Cc�?             <@0       ;                    �?`�Q��?             9@1       6                   �<@���Q��?             .@2       3                   �;@      �?             @������������������������       �                     �?4       5                 `f�D@�q�q�?             @������������������������       �                      @������������������������       �                     �?7       8                 �|Y=@���!pc�?             &@������������������������       �                      @9       :                 `f�>@�q�q�?             "@������������������������       �      �?             @������������������������       �                     @<       =                  x#J@z�G�z�?             $@������������������������       �                     @>       E                   �C@�q�q�?             @?       @                 `f�K@z�G�z�?             @������������������������       �                      @A       B                    >@�q�q�?             @������������������������       �                     �?C       D                 03�P@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     �?G       H                    �?�q�q�?             @������������������������       �                     �?������������������������       �                      @J       Q                    �? 7���B�?             ;@K       L                   @H@ �q�q�?             8@������������������������       �                     &@M       P                   @J@$�q-�?             *@N       O                 ���W@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     $@������������������������       �                     @������������������������       �                     @T       c                    �?����H�?U            �_@U       b                    �?���N8�?             E@V       _                   �B@HP�s��?             9@W       X                    �?���N8�?             5@������������������������       �                      @Y       Z                    1@�}�+r��?             3@������������������������       �                     $@[       \                    7@�����H�?             "@������������������������       �                     @]       ^                   �7@z�G�z�?             @������������������������       �                     �?������������������������       �                     @`       a                   �C@      �?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     1@d       �                    �?�IєX�?6            @U@e       h                    4@ ��Ou��?2            �S@f       g                    &@r�q��?             @������������������������       �                     �?������������������������       �                     @i       j                 �|Y=@�X�<ݺ?.             R@������������������������       �                     7@k       �                   @F@Hm_!'1�?             �H@l       q                    �?�KM�]�?             C@m       p                 hf�2@؇���X�?             @n       o                 X�l@@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @r       s                   �?@��a�n`�?             ?@������������������������       �                     "@t       {                    �?��2(&�?             6@u       z                   @D@�����H�?             2@v       y                   @A@��S�ۿ?
             .@w       x                 `fF)@      �?              @������������������������       �                     @������������������������       ��q�q�?             @������������������������       �                     @������������������������       ��q�q�?             @|       }                   �7@      �?             @������������������������       �                     �?~       �                   �:@�q�q�?             @       �                   �@@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     �?������������������������       �                     &@������������������������       �                     @�       �                    �?�x�W�?�             w@������������������������       �                     @�       �                    �?�o(���?�            �v@�       �                    �?�i#[��??             U@�       �                    �?�I� �?#             G@�       �                    �?tk~X��?             B@�       �                    �?"pc�
�?            �@@�       �                 �|Y7@      �?              @������������������������       �                     �?������������������������       �                     �?�       �                 �̌@�חF�P�?             ?@�       �                  ��@P���Q�?             4@�       �                  �[@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     1@�       �                 �� @���|���?             &@�       �                 Ь* @և���X�?             @�       �                    �?���Q��?             @������������������������       �                     �?�       �                 �?�@      �?             @������������������������       �                     �?�       �                   �8@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                      @������������������������       �                     @�       �                    $@�q�q�?             @������������������������       �                     �?������������������������       �                      @�       �                 �A7@z�G�z�?             $@�       �                 �|�:@���Q��?             @������������������������       �                     �?�       �                 �I5@      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     @�       �                    �?�d�����?             C@�       �                   �,@�û��|�?             7@������������������������       �                      @�       �                    �?�q�q�?             5@������������������������       �                     @�       �                    �?j���� �?             1@�       �                 �|�>@�q�q�?             @������������������������       �                      @������������������������       �                     �?�       �                    �?X�Cc�?
             ,@�       �                 �|�<@      �?             $@������������������������       �                     @�       �                 ���.@r�q��?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     @�       �                 ��T?@��S�ۿ?
             .@������������������������       �                      @�       �                 ��p@@؇���X�?             @������������������������       �                     �?������������������������       �                     @�       *                   �?R���Q�?�            �q@�       �                    $@Tb.��?�            @o@������������������������       �                     @�       '                0��F@&!��Ji�?�            �n@�       �                    �?\���(\�?�             n@�       �                    �?�������?             >@�       �                 �|Y=@8�Z$���?             :@�       �                    <@X�<ݚ�?             "@�       �                 �&�)@����X�?             @�       �                   �1@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @������������������������       �                      @������������������������       �                     1@�       �                   �2@      �?             @������������������������       �                     �?������������������������       �                     @�       �                    �?�̐d��?�            @j@�       �                    �?ܷ��?��?             =@�       �                 �|Y=@�LQ�1	�?             7@������������������������       �                     �?�       �                 �|Y>@�C��2(�?             6@�       �                 ��(@�����H�?             2@�       �                  s�@8�Z$���?	             *@������������������������       �                     @������������������������       �z�G�z�?             $@������������������������       �                     @������������������������       �                     @������������������������       �                     @�                           �?`����e�?v            �f@�       �                 �?�@(Q��w��?e             c@�       �                   �;@p=
ףp�?8             T@�       �                 ��@4?,R��?             B@�       �                 `f�@�q�q�?             @�       �                    6@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     �?�       �                 �1@�C��2(�?            �@@�       �                   �:@؇���X�?             5@�       �                 �?$@ףp=
�?             4@�       �                 ���@�X�<ݺ?             2@�       �                 ���@z�G�z�?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     *@�       �                   �3@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     �?������������������������       �        	             (@�       �                 ���@���7�?             F@������������������������       �                     3@�       �                   �?@HP�s��?             9@�       �                 �?$@P���Q�?             4@�       �                 �|Y>@�q�q�?             @������������������������       �      �?              @������������������������       �                     �?������������������������       �        
             1@�       �                   �@z�G�z�?             @�       �                 �&B@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @                       @3�@&��f���?-            @R@                         :@��S���?             .@������������������������       �                     @                        �?@�q�q�?             (@������������������������       �                     @                        �A@      �?              @������������������������       ��q�q�?             @������������������������       ����Q��?             @                      `�X#@�y��*�?&             M@	                      �|Y=@�:pΈ��?!             I@
                      ���"@�θ�?             :@                        �8@"pc�
�?             6@                        �3@�KM�]�?             3@                         2@      �?              @������������������������       �                     @������������������������       �                      @������������������������       �                     &@                         <@�q�q�?             @������������������������       �                      @������������������������       �                     �?                        �<@      �?             @������������������������       �                      @������������������������       �                      @                         �? �q�q�?             8@                      ��i @�nkK�?             7@                        @?@P���Q�?             4@������������������������       �                     ,@                        �@@r�q��?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     @������������������������       �                     �?������������������������       �                      @!      &                   �?h�����?             <@"      %                   5@�}�+r��?
             3@#      $                   3@z�G�z�?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     ,@������������������������       �                     "@(      )                �|�<@z�G�z�?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     >@�t�bh�h(h+K ��h-��R�(KM+KK��h[�B�        |@     �p@     �d@      f@       @      A@              @@       @       @       @      �?              �?       @                      �?     �d@     �a@     �T@     �X@      �?     @R@              M@      �?      .@      �?                      .@     �T@      9@     �T@      6@      ;@      "@      0@      "@      0@      @              �?      0@      @      *@      @       @      �?       @      �?              �?       @              @              @      @      �?      @      �?      �?              �?      �?                       @      @              @                      @      &@             �K@      *@       @             �G@      *@               @     �G@      &@      5@      $@      @              2@      $@      1@       @      "@      @      �?      @              �?      �?       @               @      �?               @      @       @              @      @      �?      @      @               @       @      @              @       @      @      �?       @               @      �?      �?              �?      �?              �?      �?                      �?      �?       @      �?                       @      :@      �?      7@      �?      &@              (@      �?       @      �?       @                      �?      $@              @                      @     �T@     �F@       @      D@       @      7@      �?      4@               @      �?      2@              $@      �?       @              @      �?      @      �?                      @      �?      @      �?                      @              1@      T@      @     @R@      @      @      �?              �?      @              Q@      @      7@             �F@      @      A@      @      @      �?      �?      �?              �?      �?              @              <@      @      "@              3@      @      0@       @      ,@      �?      @      �?      @               @      �?      @               @      �?      @      �?      �?               @      �?      �?      �?              �?      �?              �?              &@              @             �q@     �U@              @     �q@     �T@     �E@     �D@      .@      ?@      @      =@      @      ;@      �?      �?      �?                      �?      @      :@      �?      3@      �?       @               @      �?                      1@      @      @      @      @       @      @              �?       @       @      �?              �?       @      �?                       @       @                      @      �?       @      �?                       @       @       @      @       @              �?      @      �?      @                      �?      @              <@      $@      ,@      "@               @      ,@      @      @              $@      @      �?       @               @      �?              "@      @      @      @      @              �?      @      �?                      @      @              ,@      �?       @              @      �?              �?      @             �m@      E@      j@      E@              @      j@     �B@     �i@     �@@      7@      @      6@      @      @      @      @       @      �?       @               @      �?              @                       @      1@              �?      @      �?                      @      g@      :@      :@      @      4@      @              �?      4@       @      0@       @      &@       @      @               @       @      @              @              @             �c@      7@     ``@      6@     @R@      @      ?@      @      �?       @      �?      �?      �?                      �?              �?      >@      @      2@      @      2@       @      1@      �?      @      �?      @                      �?      *@              �?      �?      �?                      �?              �?      (@              E@       @      3@              7@       @      3@      �?       @      �?      �?      �?      �?              1@              @      �?      �?      �?      �?                      �?      @              M@      .@      @       @      @              @       @              @      @      @      �?       @      @       @     �I@      @     �E@      @      4@      @      2@      @      1@       @      @       @      @                       @      &@              �?       @               @      �?               @       @       @                       @      7@      �?      6@      �?      3@      �?      ,@              @      �?              �?      @              @              �?               @              ;@      �?      2@      �?      @      �?      @                      �?      ,@              "@              �?      @      �?                      @      >@        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh$hNhJ�R�[hG        hNhG        hAKhBKhCh(h+K ��h-��R�(KK��h[�C              �?�t�bhOh`hJC       ���R�hdKhehhKh(h+K ��h-��R�(KK��hJ�C       �t�bK��R�}�(hKhrMhsh(h+K ��h-��R�(KM��hz�B(<         b                    �?J�?��?�           @�@       Q                 Ь�9@J����E�?�            pp@       P                    @���-|$�?\            @c@                            @����6Z�?X            `b@                           �?�7��?            �C@                          �9@      �?             @@       
                 ��*@����X�?             @       	                   �'@���Q��?             @������������������������       �                     �?������������������������       �      �?             @������������������������       �                      @������������������������       �                     9@������������������������       �                     @       I                 �|�=@����0�?@             [@       ,                    �?��p����?:            @X@       #                    �? s�n_Y�?"             J@                           �?      �?             8@                          �0@�8��8��?             (@������������������������       �                     @                           �?r�q��?             @                           �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @       "                    �?�q�q�?             (@       !                    �?z�G�z�?             $@                          �,@�<ݚ�?             "@������������������������       �                     �?                         �|Y6@      �?              @                          �-@      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     @������������������������       �                     �?������������������������       �                      @$       +                    �?@4և���?             <@%       &                 �|Y8@ףp=
�?             4@������������������������       �                     @'       (                 ���@      �?             0@������������������������       �                     �?)       *                 pF @��S�ۿ?             .@������������������������       �                     ,@������������������������       �                     �?������������������������       �                      @-       @                    �?���Q��?            �F@.       =                    �?���Q��?             >@/       0                 �&B@���|���?             6@������������������������       �                     @1       :                    �?�d�����?             3@2       9                 pF�!@�	j*D�?             *@3       8                 @3�@X�<ݚ�?             "@4       5                   �8@      �?              @������������������������       �                      @6       7                   �;@r�q��?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @;       <                    $@r�q��?             @������������������������       �                     �?������������������������       �                     @>       ?                    1@      �?              @������������������������       �                     @������������������������       �                     @A       F                    �?���Q��?	             .@B       C                 �!@X�<ݚ�?             "@������������������������       �                     �?D       E                 �|�;@      �?              @������������������������       �                     @������������������������       �                     @G       H                 �|�0@r�q��?             @������������������������       �                     @������������������������       �                     �?J       K                   �@@"pc�
�?             &@������������������������       �                     @L       O                    �?�q�q�?             @M       N                 `f�/@���Q��?             @������������������������       �                     @������������������������       �                      @������������������������       �                     �?������������������������       �                     @R       S                    @�~i��?F            @[@������������������������       �                     @T       a                    @����?D            @Z@U       \                     @` A�c̭?@             Y@V       W                     �?�q�q�?=             X@������������������������       �        ,            @R@X       Y                    E@�nkK�?             7@������������������������       �                     5@Z       [                   �G@      �?              @������������������������       �                     �?������������������������       �                     �?]       ^                    �?      �?             @������������������������       �                     �?_       `                    @�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @c                          �?v���%��?           |@d       �                    �?�'F����?�            �w@e       �                 ��$:@$΅9>��?�            `t@f       q                     @��c+��?�            �p@g       h                 ��Y)@�h����?&             L@������������������������       �                     4@i       p                 `��,@�8��8��?             B@j       k                 �|�<@ �Cc}�?             <@������������������������       �        
             ,@l       o                   �A@d}h���?	             ,@m       n                    �?      �?             @������������������������       �                     �?������������������������       ����Q��?             @������������������������       �                      @������������������������       �                      @r       y                   �2@�����?�            `j@s       x                 pf� @�t����?	             1@t       u                   �0@X�<ݚ�?             "@������������������������       �                      @v       w                 pf�@և���X�?             @������������������������       �                     @������������������������       �                     @������������������������       �                      @z       �                    �?�^'�ë�?|            @h@{       �                   �+@h㱪��?!            �K@|       �                 ���@@3����?              K@}       ~                 ���@`2U0*��?             9@������������������������       �        	             2@       �                 �|=@؇���X�?             @������������������������       �                      @������������������������       �z�G�z�?             @������������������������       �                     =@������������������������       �                     �?�       �                 ��@hb����?[            `a@�       �                 �|Y<@�FVQ&�?            �@@�       �                 ���@"pc�
�?             &@�       �                   �9@�q�q�?             @�       �                 �&b@z�G�z�?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @������������������������       �                     6@�       �                 �|Y=@f1r��g�?F            �Z@�       �                   �3@��<D�m�?             �H@�       �                 0S5 @z�G�z�?             @�       �                 �?�@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @�       �                   �;@���7�?             F@�       �                   �:@�IєX�?             A@�       �                   �5@      �?             @@�       �                   �4@@4և���?	             ,@������������������������       �                     @�       �                 �1@ףp=
�?             $@������������������������       �                     �?������������������������       �                     "@������������������������       �        
             2@�       �                 pb@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     $@�       �                   �F@�MWl��?&            �L@�       �                   �@�c�����?$            �J@�       �                 �&B@և���X�?             @�       �                 �|Y>@      �?             @������������������������       �      �?             @������������������������       �                      @������������������������       �                     �?�       �                 ��) @�3Ea�$�?              G@�       �                 @3�@R���Q�?             D@�       �                   @C@�d�����?             3@�       �                 �|�>@��S�ۿ?
             .@������������������������       �                      @�       �                 �?�@؇���X�?             @������������������������       �                     @������������������������       ��q�q�?             @������������������������       �                     @�       �                    ?@���N8�?             5@������������������������       �                     .@�       �                   �@@r�q��?             @������������������������       �                     �?������������������������       �                     @�       �                 ��y @      �?             @������������������������       �                     �?�       �                 ���!@���Q��?             @������������������������       �                     �?�       �                 03�0@      �?             @�       �                   �?@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @�       �                 ��";@�e�,��?!            �M@�       �                   x:@r�q��?             (@������������������������       �                     @�       �                    D@      �?              @������������������������       �                     @�       �                    H@�q�q�?             @������������������������       �                      @������������������������       �                     �?�       �                     @��k=.��?            �G@�       �                   �H@"pc�
�?             F@�       �                    �?�C��2(�?            �@@������������������������       �                     (@�       �                     �?؇���X�?             5@�       �                   �B@@�0�!��?
             1@�       �                   �<@�z�G��?             $@������������������������       �                     @������������������������       �                     @������������������������       �                     @������������������������       �                     @�       �                   @>@�eP*L��?             &@������������������������       �                     �?�       �                    �?���Q��?             $@�       �                  ��@@      �?             @������������������������       �                     �?�       �                   �O@�q�q�?             @������������������������       �                      @������������������������       �                     �?�       �                    @@�q�q�?             @�       �                   �J@      �?             @������������������������       �                      @������������������������       �                      @������������������������       �                      @�       �                    ;@�q�q�?             @������������������������       �                     �?������������������������       �                      @�       �                    �?x��}�?)            �K@�       �                     �?��
ц��?	             *@�       �                   �H@�q�q�?             @������������������������       �                     @������������������������       �                      @�       �                     @����X�?             @������������������������       �                     @�       �                 �&�)@      �?             @������������������������       �                      @������������������������       �                      @�                          H@r�q��?              E@�                          �?�p ��?            �D@�       �                   �7@b�h�d.�?            �A@������������������������       �                     3@�       �                   �@@      �?             0@�       �                     �?�q�q�?             @�       �                    7@�q�q�?             @������������������������       �                     �?�       �                 ���M@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @�                           �?z�G�z�?             $@�       �                   �B@�q�q�?             @������������������������       �                     �?�       �                  x#J@���Q��?             @������������������������       �                      @�                           F@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @������������������������       �                     @������������������������       �                     �?                          @�t����?*             Q@                        �4@�g�y��?             ?@������������������������       �                     (@                         �?�S����?             3@	                         �?�q�q�?             "@
                      �̾w@���Q��?             @������������������������       �                      @������������������������       �                     @������������������������       �                     @������������������������       �                     $@                         @$G$n��?            �B@                         @X�<ݚ�?             "@������������������������       �                     @������������������������       �                     @������������������������       �                     <@�t�bh�h(h+K ��h-��R�(KMKK��h[�B0       �z@     �q@     �M@     �i@     �G@     �Z@      D@     �Z@       @     �B@       @      >@       @      @       @      @              �?       @       @               @              9@              @      C@     �Q@      =@      Q@      &@     �D@      "@      .@      �?      &@              @      �?      @      �?      �?              �?      �?                      @       @      @       @       @      @       @              �?      @      �?      @      �?      @                      �?      @              �?                       @       @      :@       @      2@              @       @      ,@      �?              �?      ,@              ,@      �?                       @      2@      ;@      (@      2@       @      ,@      @              @      ,@      @      "@      @      @      @      @       @              �?      @              @      �?              �?                      @      �?      @      �?                      @      @      @      @                      @      @      "@      @      @              �?      @      @      @                      @      �?      @              @      �?              "@       @      @              @       @      @       @      @                       @      �?              @              (@     @X@      @               @     @X@      @     @X@      �?     �W@             @R@      �?      6@              5@      �?      �?      �?                      �?       @       @              �?       @      �?       @                      �?      @             w@      T@     t@      N@     pq@     �G@     �m@      <@     �J@      @      4@             �@@      @      9@      @      ,@              &@      @      @      @              �?      @       @       @               @             @g@      9@      (@      @      @      @               @      @      @      @                      @       @             �e@      4@     �J@       @     �J@      �?      8@      �?      2@              @      �?       @              @      �?      =@                      �?     @^@      2@      ?@       @      "@       @      @       @      @      �?      @                      �?              �?      @              6@             �V@      0@      G@      @      @      �?      �?      �?      �?                      �?      @              E@       @      @@       @      ?@      �?      *@      �?      @              "@      �?              �?      "@              2@              �?      �?              �?      �?              $@              F@      *@      D@      *@      @      @      @      @      �?      @       @                      �?     �B@      "@      A@      @      ,@      @      ,@      �?       @              @      �?      @               @      �?              @      4@      �?      .@              @      �?              �?      @              @      @              �?      @       @      �?               @       @      �?       @               @      �?              �?              @              D@      3@       @      $@              @       @      @              @       @      �?       @                      �?      C@      "@      B@       @      >@      @      (@              2@      @      ,@      @      @      @              @      @              @              @              @      @              �?      @      @       @       @      �?              �?       @               @      �?              @       @       @       @               @       @               @               @      �?              �?       @              E@      *@      @      @       @      @              @       @              @       @      @               @       @               @       @             �A@      @     �A@      @      =@      @      3@              $@      @       @      @       @      �?      �?              �?      �?              �?      �?                      @       @       @      @       @      �?              @       @       @              �?       @               @      �?              @              @                      �?      H@      4@      0@      .@              (@      0@      @      @      @       @      @       @                      @      @              $@              @@      @      @      @              @      @              <@        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh$hNhJ�v}hG        hNhG        hAKhBKhCh(h+K ��h-��R�(KK��h[�C              �?�t�bhOh`hJC       ���R�hdKhehhKh(h+K ��h-��R�(KK��hJ�C       �t�bK��R�}�(hKhrM7hsh(h+K ��h-��R�(KM7��hz�BD         ~                    �?4�<����?�           @�@       k                 ��T?@ \� ���?�            �n@       f                    @�3[�s(�?e            �b@                           @~�u���?`            �a@                           �?�G�z��?             4@                           �?      �?             2@������������������������       �                     �?                        �|>@��.k���?             1@	       
                  s@և���X�?
             ,@������������������������       �                      @                           �?      �?             (@                        �|�6@      �?             @������������������������       �                     �?                        ���@�q�q�?             @������������������������       �                     �?������������������������       �                      @                          �3@      �?              @������������������������       �                     @                        �|�9@���Q��?             @������������������������       �                     @������������������������       �                      @������������������������       �                     @������������������������       �                      @       5                     @������?R            �^@       4                    �?�LQ�1	�?#             G@       )                   �2@@�0�!��?             A@                           �9@�C��2(�?             6@                          �'@      �?             @������������������������       �                      @                          �7@      �?              @������������������������       �                     �?������������������������       �                     �?!       "                 ��Y)@�X�<ݺ?             2@������������������������       �                      @#       (                   �,@ףp=
�?             $@$       %                   �B@      �?              @������������������������       �                     @&       '                    D@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @*       -                    �?�q�q�?	             (@+       ,                    D@      �?             @������������������������       �                     @������������������������       �                     �?.       3                    D@      �?              @/       2                   �7@r�q��?             @0       1                    �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @������������������������       �                      @������������������������       �        
             (@6       Q                   �*@rOP\6�?/            @S@7       L                    �?��R[s�?            �A@8       ?                  ��@l��
I��?             ;@9       >                    �?�����H�?             "@:       ;                 ��H@r�q��?             @������������������������       �                     @<       =                 �|Y>@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @@       A                   �3@b�2�tk�?             2@������������������������       �                     @B       K                 ��"@�q�q�?	             (@C       D                    �?      �?             $@������������������������       �                     �?E       F                   �9@X�<ݚ�?             "@������������������������       �                     @G       H                   �<@r�q��?             @������������������������       �                     @I       J                   �>@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                      @M       N                   �#@      �?              @������������������������       �                     @O       P                 P��%@�q�q�?             @������������������������       �                     �?������������������������       �                      @R       e                   @D@�G��l��?             E@S       ^                    �?D�n�3�?             C@T       ]                 �=/@�q�q�?             8@U       Z                    �?�n_Y�K�?             *@V       Y                 ���,@�q�q�?             "@W       X                 �|Y6@      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     @[       \                 �|�>@      �?             @������������������������       �                      @������������������������       �                      @������������������������       �                     &@_       d                 �|�<@և���X�?	             ,@`       a                    �?z�G�z�?             $@������������������������       �                     @b       c                 `f7@���Q��?             @������������������������       �                      @������������������������       �                     @������������������������       �                     @������������������������       �                     @g       h                    )@      �?              @������������������������       �                     @i       j                    �?�q�q�?             @������������������������       �                      @������������������������       �                     �?l       m                    �?heu+��?A            �W@������������������������       �        .             Q@n       y                   �8@R�}e�.�?             :@o       v                     @r�q��?             2@p       q                    �?��S�ۿ?	             .@������������������������       �                     @r       s                 ���`@�8��8��?             (@������������������������       �                     "@t       u                 ���i@�q�q�?             @������������������������       �                     �?������������������������       �                      @w       x                    %@�q�q�?             @������������������������       �                     �?������������������������       �                      @z       {                 X�l@@      �?              @������������������������       �                     @|       }                    @z�G�z�?             @������������������������       �                     @������������������������       �                     �?       �                    ,@jN�{��?           0}@�       �                     @���Q��?             >@������������������������       �                     &@�       �                    �?p�ݯ��?
             3@������������������������       �                     �?�       �                     @�q�q�?	             2@������������������������       �                     @�       �                    @$�q-�?             *@�       �                    �?z�G�z�?             @������������������������       �                     @������������������������       �                     �?������������������������       �                      @�       0                   �?��b��?
           P{@�       �                    �? �@��:�?�            �x@�       �                     �?�C��2(�?            �K@�       �                   @@@��2(&�?
             6@������������������������       �                     &@�       �                   �E@���!pc�?             &@������������������������       �                     @������������������������       �                      @�       �                    �?�FVQ&�?            �@@�       �                     @���}<S�?             7@�       �                 `��,@      �?              @������������������������       �                     �?������������������������       �                     �?�       �                 �|Y=@���N8�?             5@�       �                   @:@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     3@������������������������       �                     $@�       -                   �?<�W�V�?�            Pu@�       �                     �?zCK��?�            �t@�       �                   �<@��>4և�?'             L@�       �                    �?z�G�z�?             $@�       �                   �;@؇���X�?             @������������������������       �                     �?�       �                 `f�D@r�q��?             @������������������������       �                     @������������������������       �                     �?�       �                    7@�q�q�?             @������������������������       �                     �?������������������������       �                      @�       �                    @@8����?!             G@�       �                   �@@П[;U��?             =@�       �                 �|Y=@�����H�?             "@������������������������       �                     �?�       �                 �|Y?@      �?              @�       �                 `fF:@؇���X�?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     �?�       �                   �F@���Q��?             4@�       �                 ��I*@�����H�?             "@������������������������       �                     �?������������������������       �                      @�       �                   @=@���|���?             &@�       �                 ��:@؇���X�?             @������������������������       �                      @�       �                    J@z�G�z�?             @�       �                 `f�;@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @�       �                   @>@      �?             @������������������������       �                      @�       �                   �J@      �?              @������������������������       �                     �?������������������������       �                     �?�       �                 ��9L@�IєX�?             1@������������������������       �        	             *@�       �                 `f�N@      �?             @������������������������       �                     �?������������������������       �                     @�       $                   �?lGts��?�            0q@�       �                    �?��0 >_�?�            `o@�       �                     @��+7��?             7@������������������������       �                     @�       �                 �|Y=@�z�G��?             4@������������������������       �                     @�       �                  s�@      �?             0@������������������������       �                      @�       �                 �|Y>@؇���X�?	             ,@�       �                   @'@����X�?             @������������������������       ����Q��?             @������������������������       �                      @������������������������       �                     @�       �                   �7@@��xQ�?�            �l@�       �                     @�]0��<�?(            �N@������������������������       �                     (@�       �                   �3@@9G��?             �H@�       �                   �2@�����?             5@������������������������       �                     *@�       �                 �?�@      �?              @������������������������       �                     @�       �                 0S5 @      �?             @������������������������       �                      @������������������������       �                      @������������������������       �                     <@�       !                0��D@�-�����?`            �d@�       �                   �;@�Iy4�%�?^            `d@�       �                     @d}h���?             <@������������������������       �                     (@�       �                   �:@      �?
             0@�       �                   �8@�����H�?             "@������������������������       �                     �?������������������������       �                      @�       �                 pb@����X�?             @������������������������       �                     @������������������������       �                      @�       �                     @�:�^���?N            �`@�       �                   �G@�㙢�c�?             7@�       �                 `fF)@���y4F�?             3@������������������������       �                     @�       �                   �*@����X�?             ,@�       �                 �|�=@���|���?             &@������������������������       �                     �?�       �                    @@�z�G��?             $@������������������������       �                      @�       �                   �A@      �?              @������������������������       ��q�q�?             @�       �                   �C@z�G�z�?             @������������������������       �                     �?������������������������       �      �?             @������������������������       �                     @������������������������       �                     @�                       ���"@@4և���?=             \@�       �                 ��@��^M}�?6            @Y@������������������������       �                     A@                         �?@t�e�í�?'            �P@                      �|Y=@��Y��]�?            �D@������������������������       �                     $@                      �|�=@�g�y��?             ?@                       sW@ ��WV�?             :@������������������������       ��q�q�?             @������������������������       �                     7@������������������������       �                     @                      @3�@8�Z$���?             :@	                        �M@և���X�?             @
                        �@      �?             @������������������������       �                     �?                        @C@���Q��?             @                      �?�@      �?             @������������������������       �                     �?������������������������       ��q�q�?             @������������������������       �                     �?������������������������       �                     �?                        @F@�}�+r��?	             3@������������������������       �                     .@                        �G@      �?             @������������������������       �                     �?������������������������       �                     @                      �|�=@���!pc�?             &@                      ���(@      �?              @                        �<@z�G�z�?             @������������������������       �                      @                      �|Y=@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     @                         �?@�q�q�?             @������������������������       �                      @������������������������       �                     �?"      #                �|�;@      �?             @������������������������       �                      @������������������������       �                      @%      &                �|�>@�8��8��?             8@������������������������       �        	             ,@'      ,                    @z�G�z�?             $@(      )                  �7@�<ݚ�?             "@������������������������       �                      @*      +                  �@@����X�?             @������������������������       �                      @������������������������       �                     @������������������������       �                     �?.      /                  �G@z�G�z�?             $@������������������������       �                      @������������������������       �                      @1      6                  �6@������?            �D@2      3                   �?      �?             @������������������������       �                     �?4      5                   3@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                    �B@�t�bh�h(h+K ��h-��R�(KM7KK��h[�Bp        |@     �p@      N@      g@     �J@     �X@      G@     @X@      &@      "@      "@      "@              �?      "@       @      @       @               @      @      @      �?      @              �?      �?       @      �?                       @      @      @      @               @      @              @       @              @               @             �A@      V@      @      D@      @      <@       @      4@      �?      @               @      �?      �?              �?      �?              �?      1@               @      �?      "@      �?      @              @      �?      �?      �?                      �?               @      @       @      �?      @              @      �?              @      @      �?      @      �?      �?              �?      �?                      @       @                      (@      =@      H@      "@      :@       @      3@      �?       @      �?      @              @      �?       @               @      �?                      @      @      &@              @      @      @      @      @      �?              @      @      @              �?      @              @      �?       @      �?                       @       @              �?      @              @      �?       @      �?                       @      4@      6@      0@      6@       @      0@       @      @      @      @      �?      @              @      �?              @               @       @               @       @                      &@       @      @       @       @      @              @       @               @      @                      @      @              @      �?      @               @      �?       @                      �?      @     �U@              Q@      @      3@      @      .@      �?      ,@              @      �?      &@              "@      �?       @      �?                       @       @      �?              �?       @              @      @      @              �?      @              @      �?             @x@     �S@      (@      2@              &@      (@      @              �?      (@      @              @      (@      �?      @      �?      @                      �?       @             �w@     �N@     u@     �M@      I@      @      3@      @      &@               @      @              @       @              ?@       @      5@       @      �?      �?              �?      �?              4@      �?      �?      �?      �?                      �?      3@              $@             �q@      K@     pq@      J@      A@      6@       @       @      �?      @              �?      �?      @              @      �?              �?       @      �?                       @      @@      ,@      0@      *@       @      �?      �?              @      �?      @      �?      @                      �?      �?               @      (@      �?       @      �?                       @      @      @      @      �?       @              @      �?      �?      �?              �?      �?              @              �?      @               @      �?      �?              �?      �?              0@      �?      *@              @      �?              �?      @             �n@      >@     �k@      <@      1@      @      @              ,@      @              @      ,@       @       @              (@       @      @       @      @       @       @              @             �i@      6@     �M@       @      (@             �G@       @      3@       @      *@              @       @      @               @       @               @       @              <@             `b@      4@      b@      2@      6@      @      (@              $@      @       @      �?              �?       @               @      @              @       @             �^@      (@      3@      @      .@      @      @              $@      @      @      @              �?      @      @       @              @      @      �?       @      @      �?      �?              @      �?      @              @              Z@       @      X@      @      A@              O@      @      D@      �?      $@              >@      �?      9@      �?       @      �?      7@              @              6@      @      @      @      @      @              �?      @       @      @      �?      �?               @      �?              �?      �?              2@      �?      .@              @      �?              �?      @               @      @      @      �?      @      �?       @               @      �?              �?       @              @              �?       @               @      �?               @       @               @       @              6@       @      ,@               @       @      @       @       @              @       @               @      @              �?               @       @       @                       @     �C@       @       @       @              �?       @      �?       @                      �?     �B@        �t�bub��     hhubh)��}�(hhhhhNhKhKhG        hh$hNhJg}�XhG        hNhG        hAKhBKhCh(h+K ��h-��R�(KK��h[�C              �?�t�bhOh`hJC       ���R�hdKhehhKh(h+K ��h-��R�(KK��hJ�C       �t�bK��R�}�(hKhrM3hsh(h+K ��h-��R�(KM3��hz�B(C         �                     @^IB�A��?�           @�@       }                    �?�/����?�            `t@                         ��[+@��0u���?�             n@                           �?v���EO�?-            �Q@                        ��Y)@�<ݚ�?             2@                          �J@�����H�?             "@������������������������       �                      @������������������������       �                     �?	       
                   �B@�q�q�?             "@������������������������       �                     @                           D@      �?             @������������������������       �                     @������������������������       �                     �?                           5@ �h�7W�?!            �J@                           &@z�G�z�?             @                          �1@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @                          @A@ �q�q�?             H@                            �?@4և���?             <@������������������������       �                     @                          �@@HP�s��?             9@                        �|Y=@���N8�?             5@������������������������       �                      @                        �|�=@$�q-�?             *@                           @z�G�z�?             @������������������������       �                     @������������������������       �                     �?������������������������       �                      @������������������������       �      �?             @������������������������       �                     4@!       f                     �?V1���?p             e@"       Q                   @F@�4�����?V             _@#       8                    �?R�}e�.�?7            �S@$       7                    �?z�G�z�?             >@%       6                  "�`@��+7��?             7@&       3                 �DhF@��s����?             5@'       (                 0C�;@�q�q�?             "@������������������������       �                     @)       *                   �<@      �?             @������������������������       �                     �?+       ,                 �|�;@���Q��?             @������������������������       �                     �?-       .                  �>@      �?             @������������������������       �                     �?/       0                    �?�q�q�?             @������������������������       �                     �?1       2                   �A@      �?              @������������������������       �                     �?������������������������       �                     �?4       5                    �?�8��8��?	             (@������������������������       �                     &@������������������������       �                     �?������������������������       �                      @������������������������       �                     @9       :                    �?     ��?!             H@������������������������       �                     0@;       >                 `fF<@     ��?             @@<       =                 03:@$�q-�?             *@������������������������       �                     �?������������������������       �                     (@?       B                  x#J@�d�����?             3@@       A                   �;@�����H�?             "@������������������������       �                     �?������������������������       �                      @C       J                 03�P@���Q��?             $@D       E                    9@���Q��?             @������������������������       �                     �?F       G                    A@      �?             @������������������������       �                      @H       I                 `�iJ@      �?              @������������������������       �                     �?������������������������       �                     �?K       L                    �?z�G�z�?             @������������������������       �                     �?M       N                 03U@      �?             @������������������������       �                      @O       P                    �?      �?              @������������������������       �                     �?������������������������       �                     �?R       S                    �?��c:�?             G@������������������������       �        
             0@T       _                    �?d��0u��?             >@U       ^                 @�pX@��
ц��?             *@V       W                   �G@�q�q�?             "@������������������������       �                     �?X       ]                    �?      �?              @Y       \                   �O@      �?             @Z       [                  ��@@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     �?������������������������       �                     @������������������������       �                     @`       a                   �G@�t����?             1@������������������������       �                     $@b       c                   @>@����X�?             @������������������������       �                     @d       e                   @J@�q�q�?             @������������������������       �                     �?������������������������       �                      @g       x                   �:@��S���?            �F@h       s                    �?���@M^�?             ?@i       n                    5@�q�q�?	             (@j       m                 ���.@և���X�?             @k       l                 ���,@      �?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     @o       p                   �1@z�G�z�?             @������������������������       �                      @q       r                    �?�q�q�?             @������������������������       �                     �?������������������������       �                      @t       w                   �6@�d�����?	             3@u       v                 ��m1@      �?              @������������������������       �                     @������������������������       �                     @������������������������       �                     &@y       z                 0S�<@؇���X�?             ,@������������������������       �                     @{       |                    0@      �?              @������������������������       �                      @������������������������       �                     @~       �                    �?��T|n�?6            �U@       �                    �?      �?             H@������������������������       �                    �@@�       �                     �?z�G�z�?             .@�       �                 м{L@z�G�z�?             $@������������������������       �                     �?�       �                 pU�t@�����H�?             "@������������������������       �                      @������������������������       �                     �?�       �                    0@z�G�z�?             @������������������������       �                     �?������������������������       �                     @�       �                     �?�˹�m��?             C@������������������������       �        
             2@�       �                    �?R���Q�?             4@������������������������       �        	             .@�       �                    *@���Q��?             @������������������������       �                      @������������������������       �                     @�       �                 pff@�%����?�             x@�       �                    �?�����?(            �O@�       �                 ���@      �?             8@�       �                 03S@     ��?	             0@������������������������       �                     @�       �                 �|�9@�θ�?             *@������������������������       �                      @�       �                    �?�C��2(�?             &@������������������������       �                     �?������������������������       �                     $@������������������������       �                      @�       �                 �|Y;@$�q-�?            �C@�       �                  ��	@�S����?             3@�       �                    6@      �?             @������������������������       �                      @������������������������       �                      @�       �                    �?��S�ۿ?             .@������������������������       �                      @�       �                    �?$�q-�?             *@�       �                   �5@�����H�?             "@������������������������       �                     @�       �                   �7@      �?             @�       �                    �?�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     �?������������������������       �                     @������������������������       �                     4@�       $                @3�4@P�J>_�?�            0t@�       �                    @��i,��?�            @p@�       �                    �?$�q-�?             *@������������������������       �                     @�       �                    @r�q��?             @������������������������       �                     �?������������������������       �                     @�       �                    �?�@U����?�            �n@�       �                    �?���Q��?,            �R@�       �                 0C�3@      �?             H@�       �                 �|�=@��<b���?             G@�       �                    �?,���i�?            �D@�       �                    �?�X�<ݺ?             B@�       �                    �? >�֕�?            �A@������������������������       �                     8@�       �                 @q"@"pc�
�?             &@�       �                 P�@ףp=
�?             $@������������������������       �                     @�       �                   �8@r�q��?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     �?������������������������       �                     �?�       �                 �|�:@���Q��?             @������������������������       �                      @������������������������       �                     @������������������������       �                     @������������������������       �                      @�       �                 �|�<@�q�q�?             ;@�       �                    4@r�q��?             (@�       �                    �?����X�?             @�       �                    '@r�q��?             @������������������������       �                     @�       �                 �&�)@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     �?������������������������       �                     @�       �                    �?��S���?	             .@������������������������       �                     @�       �                   �D@�q�q�?             (@�       �                 �|Y>@�<ݚ�?             "@������������������������       �                     @�       �                    A@���Q��?             @�       �                 03C3@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                      @������������������������       �                     @�       #                   �?x�g���?s            �e@�       �                 �?�@Ԫ2��?r            `e@�       �                    �?     �?+             P@�       �                    �?���N8�?*            �O@������������������������       �                      @�       �                 �1@�.ߴ#�?(            �N@�       �                   �:@l��\��?             A@������������������������       �                     $@�       �                    �?      �?             8@�       �                  s�@�IєX�?
             1@������������������������       �                     @�       �                 X��A@�C��2(�?             &@������������������������       �ףp=
�?             $@������������������������       �                     �?�       �                 ��@����X�?             @������������������������       �                      @�       �                 �|Y?@���Q��?             @�       �                   �;@�q�q�?             @������������������������       �                     �?�       �                 �|�<@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @������������������������       �                     ;@������������������������       �                     �?�       �                    �?�!�z�0�?G            �Z@�       �                 03�-@և���X�?             @������������������������       �                      @�       �                 ؼC1@z�G�z�?             @������������������������       �                     @�       �                   �2@      �?              @������������������������       �                     �?������������������������       �                     �?�                           �?Ș����?B             Y@������������������������       �                     @      "                   D@r�q��??             X@                      ���!@�Y�����?6            �T@                         C@�\�u��?            �I@                      ��) @������?            �F@                      @3�@x�����?            �C@                        �=@����X�?             ,@������������������������       �                     @      	                  �?@���Q��?             $@������������������������       �                     @
                         �?؇���X�?             @������������������������       �      �?             @������������������������       �                     @                        �4@�J�4�?             9@                        �1@�q�q�?             @������������������������       �                     �?������������������������       �                      @                        @?@�C��2(�?             6@������������������������       �                     0@                        �@@�q�q�?             @������������������������       �                      @������������������������       �                     @                         8@�q�q�?             @������������������������       �                      @������������������������       �                     @������������������������       ��q�q�?             @      !                   �?      �?             @@                        �<@�IєX�?             1@������������������������       �        
             *@                       �|Y=@      �?             @                      ���"@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @������������������������       �        
             .@������������������������       �        	             *@������������������������       �                     �?%      2                   @�����?&            �O@&      -                   �?�q�q�?
             2@'      *                   @����X�?             @(      )                   @      �?              @������������������������       �                     �?������������������������       �                     �?+      ,                   @z�G�z�?             @������������������������       �                     �?������������������������       �                     @.      /                   @�C��2(�?             &@������������������������       �                      @0      1                �̤=@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                    �F@�t�bh�h(h+K ��h-��R�(KM3KK��h[�B0       �z@     �q@     �`@      h@     �]@     �^@      K@      1@      @      ,@      �?       @               @      �?              @      @              @      @      �?      @                      �?      I@      @      @      �?      �?      �?      �?                      �?      @              G@       @      :@       @      @              7@       @      4@      �?       @              (@      �?      @      �?      @                      �?       @              @      �?      4@              P@     @Z@      D@      U@      5@     �L@      @      8@      @      1@      @      1@      @      @              @      @      @      �?               @      @              �?       @       @      �?              �?       @              �?      �?      �?              �?      �?              �?      &@              &@      �?               @                      @      .@     �@@              0@      .@      1@      �?      (@      �?                      (@      ,@      @       @      �?              �?       @              @      @       @      @      �?              �?      @               @      �?      �?              �?      �?              @      �?      �?              @      �?       @              �?      �?      �?                      �?      3@      ;@              0@      3@      &@      @      @      @      @      �?               @      @       @       @      �?       @      �?                       @      �?                      @      @              (@      @      $@               @      @              @       @      �?              �?       @              8@      5@      (@      3@      @      @      @      @      @      �?              �?      @                      @      @      �?       @               @      �?              �?       @              @      ,@      @      @              @      @                      &@      (@       @      @              @       @               @      @              .@     �Q@      (@      B@             �@@      (@      @       @       @              �?       @      �?       @                      �?      @      �?              �?      @              @     �A@              2@      @      1@              .@      @       @               @      @             @r@     �W@     �L@      @      5@      @      *@      @      @              $@      @               @      $@      �?              �?      $@               @              B@      @      0@      @       @       @       @                       @      ,@      �?       @              (@      �?       @      �?      @              @      �?       @      �?              �?       @              �?              @              4@             `m@      V@     @f@     �T@      �?      (@              @      �?      @      �?                      @      f@     �Q@      >@     �F@      (@      B@      $@      B@      @      B@       @      A@       @     �@@              8@       @      "@      �?      "@              @      �?      @      �?                      @      �?                      �?      @       @               @      @              @               @              2@      "@      $@       @      @       @      @      �?      @               @      �?              �?       @                      �?      @               @      @      @              @      @       @      @              @       @      @       @      �?       @                      �?               @      @             `b@      9@     `b@      8@     �N@      @      N@      @       @              M@      @      ?@      @      $@              5@      @      0@      �?      @              $@      �?      "@      �?      �?              @       @       @              @       @      �?       @              �?      �?      �?      �?                      �?       @              ;@              �?             �U@      5@      @      @       @              �?      @              @      �?      �?      �?                      �?     �T@      1@      @             �S@      1@     �P@      1@     �A@      0@     �@@      (@      ?@       @      $@      @      @              @      @              @      @      �?      @      �?      @              5@      @      �?       @      �?                       @      4@       @      0@              @       @               @      @               @      @       @                      @       @      @      ?@      �?      0@      �?      *@              @      �?      �?      �?      �?                      �?       @              .@              *@                      �?     �L@      @      (@      @       @      @      �?      �?      �?                      �?      �?      @      �?                      @      $@      �?       @               @      �?       @                      �?     �F@        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh$hNhJ	�tlhG        hNhG        hAKhBKhCh(h+K ��h-��R�(KK��h[�C              �?�t�bhOh`hJC       ���R�hdKhehhKh(h+K ��h-��R�(KK��hJ�C       �t�bK��R�}�(hKhrM;hsh(h+K ��h-��R�(KM;��hz�B�D         �                    �?F�`�E��?�           @�@       3                     �?���)��?S           ��@                           �?     .�?J             `@������������������������       �                    �I@       .                   �J@\I�~�?+            @S@                           �?������?%            �O@       
                    �?r�q��?             (@       	                    C@      �?              @������������������������       �                     @������������������������       �                     �?                          �H@      �?             @������������������������       �                     �?������������������������       �                     @                        03:@�~8�e�?            �I@������������������������       �                     @       -                   �G@nM`����?             G@       ,                   �F@)O���?             B@                           �?     ��?             @@                        �|�?@���N8�?             5@                          �<@�n_Y�K�?             *@                          �;@؇���X�?             @������������������������       �                     @                        `f�D@      �?             @������������������������       �                     @������������������������       �                     �?                        �|Y=@�q�q�?             @������������������������       �                      @                        `f�>@      �?             @������������������������       �                      @������������������������       �                      @������������������������       �                      @        %                 `�iJ@���!pc�?             &@!       "                   @B@      �?             @������������������������       �                     �?#       $                  x#J@�q�q�?             @������������������������       �                     �?������������������������       �                      @&       '                    7@؇���X�?             @������������������������       �                     @(       +                 ���M@      �?             @)       *                    @@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @������������������������       �                     @������������������������       �                     $@/       0                   @A@@4և���?             ,@������������������������       �                     (@1       2                   �O@      �?              @������������������������       �                     �?������������������������       �                     �?4       _                     @�����?	           �y@5       Z                   @B@&S��:�?B             Y@6       Y                    �?���=A�?3             S@7       <                    �?F�����?2            @R@8       9                 0S�<@      �?              @������������������������       �                     @:       ;                    �?      �?              @������������������������       �                     �?������������������������       �                     �?=       @                    6@�7�֥��?,            @P@>       ?                    �?      �?	             0@������������������������       �                      @������������������������       �                      @A       D                    :@�J��%�?#            �H@B       C                    �?ףp=
�?             $@������������������������       �      �?              @������������������������       �                      @E       V                   �7@�n_Y�K�?            �C@F       I                   �(@:ɨ��?            �@@G       H                    �?؇���X�?
             ,@������������������������       �                      @������������������������       �                     (@J       K                 �|�<@D�n�3�?             3@������������������������       �                     @L       M                    �?      �?
             0@������������������������       �                     @N       U                    1@z�G�z�?             $@O       P                 �|�=@����X�?             @������������������������       �                     �?Q       T                   @@@r�q��?             @R       S                   �>@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @������������������������       �                     @W       X                    �?r�q��?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     @[       ^                    �?�8��8��?             8@\       ]                    L@���Q��?             @������������������������       �                      @������������������������       �                     @������������������������       �                     3@`       �                 �T)D@t�n_Y��?�            �s@a       b                 03�@&ӴO���?�            �r@������������������������       �                     8@c       v                   �3@@�H�-��?�            pq@d       k                    �?��.k���?             A@e       h                    �?8�Z$���?	             *@f       g                 �&�)@      �?             @������������������������       �                     @������������������������       �                     �?i       j                 ��y.@�����H�?             "@������������������������       �                      @������������������������       �                     �?l       q                 0S5 @�q�q�?             5@m       n                 �?�@X�<ݚ�?             "@������������������������       �                     @o       p                    1@r�q��?             @������������������������       �      �?              @������������������������       �                     @r       s                    �?r�q��?             (@������������������������       �                     "@t       u                    �?�q�q�?             @������������������������       �                      @������������������������       �                     �?w       �                    �?�]?��?�            �n@x                        �̌@`��}3��?#            �J@y       ~                 �|>@�����H�?             ;@z       {                    �?`2U0*��?             9@������������������������       �                     2@|       }                 �|�;@؇���X�?             @������������������������       �                     @������������������������       �                     �?������������������������       �                      @�       �                    �?��
ц��?             :@������������������������       �                      @�       �                 `�X!@      �?             8@�       �                 @3�@z�G�z�?             $@�       �                 �?�@      �?             @������������������������       �                     �?�       �                   �8@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     @�       �                 �|�;@����X�?             ,@������������������������       �                     @�       �                    �?�C��2(�?             &@������������������������       �                      @�       �                   �D@�����H�?             "@������������������������       �                      @������������������������       �                     �?�       �                   �>@�8��8��?{             h@�       �                    �?�8��8��?]             b@�       �                   �<@P�R�`M�?S            ``@�       �                 ��q1@��S�ۿ?&             N@�       �                 �1@�}�+r��?$            �L@�       �                   �5@R���Q�?             4@�       �                    �?�q�q�?             @������������������������       �                      @�       �                 �?$@      �?             @������������������������       �                      @������������������������       �                      @�       �                   �:@@4և���?
             ,@������������������������       �                     "@�       �                   �;@z�G�z�?             @������������������������       �                     �?������������������������       �                     @������������������������       �                    �B@�       �                   �4@�q�q�?             @������������������������       �                     �?������������������������       �                      @�       �                 �|Y=@�Z��L��?-            �Q@�       �                 ���@      �?             @������������������������       �                     �?������������������������       �                     @�       �                    �?pH����?*            �P@�       �                 �|�=@�L���?            �B@�       �                    �?�8��8��?             B@�       �                 ���@�r����?             .@������������������������       �                     @�       �                   @@      �?              @������������������������       ����Q��?             @������������������������       �                     @�       �                 ��(@���N8�?             5@�       �                 03�@�IєX�?	             1@������������������������       �                      @������������������������       ���S�ۿ?             .@������������������������       �                     @������������������������       �                     �?�       �                 ��) @�r����?             >@�       �                  sW@`2U0*��?             9@�       �                 �|�=@�q�q�?             @�       �                 ��@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     �?������������������������       �                     6@�       �                 �|�=@���Q��?             @�       �                 �̜!@      �?             @������������������������       �                      @������������������������       �                      @������������������������       �                     �?������������������������       �        
             *@�       �                    �?r�qG�?             H@�       �                 �?�@��i#[�?             E@�       �                 �&B@�IєX�?             1@������������������������       �                     (@�       �                   �@z�G�z�?             @������������������������       �                     �?������������������������       �                     @�       �                 @3�@�q�����?             9@�       �                   �?@r�q��?             (@������������������������       �                     @�       �                   �D@�q�q�?             @�       �                   �A@���Q��?             @������������������������       �      �?              @������������������������       ��q�q�?             @������������������������       �                     �?�       �                 pf� @8�Z$���?             *@�       �                   @F@"pc�
�?             &@������������������������       �                     @�       �                   �G@���Q��?             @������������������������       �                      @������������������������       �                     @������������������������       �                      @������������������������       �                     @�       �                 �|�<@�����H�?             "@�       �                    ;@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @�                           @�����?n            �e@�       �                   �8@������?:            �V@�       �                    �? qP��B�?            �E@�       �                    �?�}�+r��?             3@�       �                 ��c@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     0@������������������������       �                     8@�       �                    �?z�J��?            �G@�       �                    �?��Q��?             4@������������������������       �                     @�       �                    �?@4և���?             ,@�       �                 @�ys@�����H�?             "@������������������������       �                      @������������������������       �                     �?������������������������       �                     @�                          P@��}*_��?             ;@�                          �<@$��m��?             :@�       �                    �?�eP*L��?             &@�       �                   �A@      �?             @������������������������       �                     @������������������������       �                     �?�       �                   �8@����X�?             @������������������������       �                     �?�       �                    �?r�q��?             @�       �                   �B@z�G�z�?             @�       �                    �?�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                      @������������������������       �                     �?      
                   �?z�G�z�?             .@                      0�:P@"pc�
�?	             &@������������������������       �                     @                        @D@�q�q�?             @������������������������       �                     �?                        �J@z�G�z�?             @������������������������       �                     @      	                   �?      �?              @������������������������       �                     �?������������������������       �                     �?                      ���`@      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     �?      "                   @�A����?4            �T@                         �?
j*D>�?             :@                         �?��.k���?             1@                      ��*4@���|���?             &@                         �?      �?              @������������������������       �                     @                         �?z�G�z�?             @                        �&@      �?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     �?������������������������       �                     @                         �?r�q��?             @������������������������       �                     @                          @�q�q�?             @������������������������       �                     �?������������������������       �                      @       !                   @�<ݚ�?             "@������������������������       �                      @������������������������       �                     @#      2                ��.@؇���X�?%             L@$      +                   �?      �?
             ,@%      &                   �?�q�q�?             @������������������������       �                     @'      (                   �?�q�q�?             @������������������������       �                     �?)      *                   �?      �?              @������������������������       �                     �?������������������������       �                     �?,      /                   �?      �?              @-      .                ��y&@z�G�z�?             @������������������������       �                     �?������������������������       �                     @0      1                   @�q�q�?             @������������������������       �                      @������������������������       �                     �?3      :                ���4@�Ń��̧?             E@4      9                   �?z�G�z�?             @5      6                   �?�q�q�?             @������������������������       �                     �?7      8                032@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @������������������������       �                    �B@�t�bh�h(h+K ��h-��R�(KM;KK��h[�B�       �z@     �q@     pu@     �h@     �F@     �T@             �I@     �F@      @@      @@      ?@      $@       @      @      �?      @                      �?      @      �?              �?      @              6@      =@      @              1@      =@      1@      3@      *@      3@      @      0@      @       @      �?      @              @      �?      @              @      �?              @       @       @               @       @               @       @                       @       @      @       @       @      �?              �?       @      �?                       @      @      �?      @              @      �?      �?      �?              �?      �?               @              @                      $@      *@      �?      (@              �?      �?              �?      �?             �r@     �\@     @R@      ;@     �I@      9@      H@      9@      @      �?      @              �?      �?              �?      �?             �D@      8@       @       @               @       @             �@@      0@      "@      �?      �?      �?       @              8@      .@      7@      $@      (@       @               @      (@              &@       @      @               @       @              @       @       @      @       @              �?      @      �?       @      �?       @                      �?      @              @              �?      @      �?                      @      @              6@       @      @       @               @      @              3@              l@     �U@      l@     �S@      8@              i@     �S@      0@      2@       @      &@      �?      @              @      �?              �?       @               @      �?              ,@      @      @      @      @              �?      @      �?      �?              @      $@       @      "@              �?       @               @      �?              g@     �N@      1@      B@      @      8@      �?      8@              2@      �?      @              @      �?               @              ,@      (@       @              (@      (@       @       @       @       @      �?              �?       @      �?                       @      @              @      $@      @              �?      $@               @      �?       @               @      �?             �d@      9@     �`@      (@     �]@      (@      L@      @      K@      @      1@      @      @       @       @               @       @       @                       @      *@      �?      "@              @      �?              �?      @             �B@               @      �?              �?       @             �O@       @      @      �?              �?      @              N@      @      A@      @     �@@      @      *@       @      @              @       @      @       @      @              4@      �?      0@      �?       @              ,@      �?      @              �?              :@      @      8@      �?       @      �?      �?      �?      �?                      �?      �?              6@               @      @       @       @               @       @                      �?      *@             �A@      *@      =@      *@      0@      �?      (@              @      �?              �?      @              *@      (@       @      $@              @       @      @       @      @      �?      �?      �?       @              �?      &@       @      "@       @      @              @       @               @      @               @              @              �?       @      �?       @               @      �?                      @     �T@     @V@      8@     �P@      �?      E@      �?      2@      �?       @               @      �?                      0@              8@      7@      8@      *@      @              @      *@      �?       @      �?       @                      �?      @              $@      1@      "@      1@      @      @      �?      @              @      �?              @       @              �?      @      �?      @      �?       @      �?              �?       @               @              �?              @      (@       @      "@              @       @      @      �?              �?      @              @      �?      �?              �?      �?              �?      @              @      �?              �?             �M@      7@      &@      .@      "@       @      @      @      �?      @              @      �?      @      �?      @      �?                      @              �?      @              @      �?      @               @      �?              �?       @               @      @       @                      @      H@       @      @      @      @       @      @              �?       @              �?      �?      �?              �?      �?              @      @      �?      @      �?                      @       @      �?       @                      �?     �D@      �?      @      �?       @      �?      �?              �?      �?      �?                      �?       @             �B@        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh$hNhJ�ޡhG        hNhG        hAKhBKhCh(h+K ��h-��R�(KK��h[�C              �?�t�bhOh`hJC       ���R�hdKhehhKh(h+K ��h-��R�(KK��hJ�C       �t�bK��R�}�(hKhrMOhsh(h+K ��h-��R�(KMO��hz�BHI                           �R@�SF�o��?�           @�@       c                    �?�CV�m�?�           ��@       P                   �B@6�B�w�?�            @i@       I                 м�9@p����?u            �e@       .                    �?�b��-8�?W            �_@       -                   �>@�3Ea�$�?=             W@       ,                 03�7@�?a/��?7            �T@       	                  �[@"�W1��?6            �T@������������������������       �                     @
                        ���@�A+K&:�?2             S@������������������������       �                      @       )                   @,@x!'ǯ�?1            �R@       $                 ��&@"pc�
�?+            �P@       #                 �|�=@��[�8��?             �I@                            @r�q��?             H@������������������������       �                     @       "                 �|�<@:	��ʵ�?            �F@                           !@l��
I��?             ;@������������������������       �                     �?                           �?R�}e�.�?             :@������������������������       �                     "@       !                 �[$@j���� �?	             1@                         @�"@      �?             0@                           5@��
ц��?             *@������������������������       �                     @                        �?�@�z�G��?             $@                          �7@���Q��?             @������������������������       �                     @������������������������       �                      @                           9@z�G�z�?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     @������������������������       �                     �?������������������������       �                     2@������������������������       �                     @%       &                   �7@��S�ۿ?             .@������������������������       �                      @'       (                   �9@؇���X�?             @������������������������       �      �?              @������������������������       �                     @*       +                 ���.@      �?              @������������������������       �                     @������������������������       �                     @������������������������       �                     �?������������������������       �                     "@/       F                    @��.k���?             A@0       1                    @*;L]n�?             >@������������������������       �                     @2       =                   �;@|��?���?             ;@3       <                    �?���!pc�?             &@4       5                     @�z�G��?             $@������������������������       �                     �?6       ;                 03�-@�q�q�?             "@7       8                 H�N&@���Q��?             @������������������������       �                     �?9       :                   �-@      �?             @������������������������       �                      @������������������������       �                      @������������������������       �                     @������������������������       �                     �?>       A                 �|�=@     ��?             0@?       @                 pF�-@      �?             (@������������������������       �                     @������������������������       �                     "@B       C                    �?      �?             @������������������������       �                     �?D       E                 `fV6@�q�q�?             @������������������������       �                      @������������������������       �                     �?G       H                    �?      �?             @������������������������       �                     @������������������������       �                     �?J       K                    �?���}<S�?             G@������������������������       �                    �C@L       O                    @և���X�?             @M       N                 ��T?@      �?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     @Q       b                     @��S���?             >@R       W                   �*@���!pc�?             6@S       T                   �'@�q�q�?             @������������������������       �                      @U       V                    D@      �?             @������������������������       �                      @������������������������       �                      @X       [                    �?      �?	             0@Y       Z                   �H@�8��8��?             (@������������������������       �                     &@������������������������       �                     �?\       a                    �?      �?             @]       `                    �?�q�q�?             @^       _                 ��yD@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     �?������������������������       �                     �?������������������������       �                      @d       o                    ,@�W��?           �z@e       f                     @�5��?             ;@������������������������       �                     @g       h                 ���4@�G��l��?             5@������������������������       �                     "@i       n                    @�8��8��?
             (@j       k                    @r�q��?             @������������������������       �                      @l       m                    @      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     @p       �                 �?�@�S� �?           �x@q       r                     @�S(��d�?\            @c@������������������������       �                     $@s       v                 ��@�8��8��?W             b@t       u                 �|Y<@"pc�
�?             &@������������������������       �                      @������������������������       �                     "@w       �                    �?`�bV��?P            �`@x       �                    �?���V��?            �F@y       �                 03s@�T|n�q�?            �E@z       �                 �|Y=@8�Z$���?            �C@{       �                  ��@X�<ݚ�?             "@|                           �?�q�q�?             @}       ~                   �6@      �?             @������������������������       �                      @������������������������       �                      @������������������������       �                      @������������������������       �                     @�       �                    �?(;L]n�?             >@�       �                 ���@@4և���?             ,@������������������������       �                     $@�       �                 �|�=@      �?             @������������������������       ��q�q�?             @������������������������       �                     �?������������������������       �                     0@�       �                 �|Y=@      �?             @������������������������       �                     �?������������������������       �                     @������������������������       �                      @�       �                    �?�zvܰ?4             V@�       �                 �?$@P��BNֱ?2            �T@������������������������       �                     H@�       �                 ��L@�#-���?            �A@�       �                   �;@�q�q�?             @������������������������       �                      @������������������������       �                     �?�       �                 �|�>@      �?             @@������������������������       �                     =@�       �                   �@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     @�       �                 @3�@ �y63��?�            �n@�       �                   �:@X�<ݚ�?             "@������������������������       �                     @�       �                   �A@�q�q�?             @������������������������       �      �?             @������������������������       �                      @�       �                     �?�2~,��?�            �m@�       �                   �<@"Ae���?#            �G@�       �                   �6@      �?              @������������������������       �                      @�       �                    �?r�q��?             @������������������������       �                      @�       �                 `f�D@      �?             @������������������������       �                     @������������������������       �                     �?�       �                    �?�(�Tw��?            �C@�       �                 03k:@     ��?             @@�       �                 X�,@@      �?             @������������������������       �                     �?������������������������       �                     @�       �                   `E@      �?             <@�       �                   �A@8����?             7@�       �                 �TA@@���!pc�?             6@�       �                   �J@�q�q�?             2@�       �                    �?և���X�?             ,@�       �                 X�lA@      �?             @������������������������       �                     @������������������������       �                     �?�       �                   `G@      �?             $@�       �                 `f�;@����X�?             @�       �                 X��B@�q�q�?             @������������������������       �      �?             @������������������������       �      �?              @������������������������       �                     �?������������������������       �                     @������������������������       �                     @������������������������       �                     @������������������������       �                     �?������������������������       �                     @�       �                 03�M@؇���X�?             @�       �                    A@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     @�                       ��.@؇���X�?|            �g@�       �                    �?F�t�K��?L            �\@�       �                 P�J.@���|���?             &@�       �                 �|Y<@      �?              @������������������������       �                     @�       �                 X�l@@�q�q�?             @�       �                 03�&@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     �?������������������������       �                     @�                          �*@6�"W�u�?E            �Y@�       �                    �?��܂O�?>            �V@�       �                 ��Y)@��f��?<            @V@�       �                   �3@�x
�2�?1            �R@�       �                 ��Y @���Q��?             $@������������������������       �                     @�       �                    $@؇���X�?             @������������������������       �                     @�       �                    &@      �?              @������������������������       �                     �?������������������������       �                     �?�       �                     @     ��?*             P@������������������������       �        	             ,@�       �                 �|�=@�:pΈ��?!             I@�       �                   �:@�X�<ݺ?             B@������������������������       �        
             3@�       �                 pf� @�t����?             1@������������������������       �                     (@�       �                 �|Y=@���Q��?             @�       �                 0S%"@�q�q�?             @������������������������       �                     �?�       �                 ���"@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @�       �                   �@@X�Cc�?             ,@�       �                 ���!@և���X�?             @�       �                 ��i @���Q��?             @�       �                    ?@      �?             @������������������������       �                      @������������������������       �                      @������������������������       �                     �?������������������������       �                      @�       �                   @F@؇���X�?             @������������������������       �                     @�       �                    G@�q�q�?             @������������������������       �                     �?������������������������       �                      @�       �                 �|�:@��S���?             .@������������������������       �                     @�       �                   @@@�q�q�?             (@������������������������       �                     @�       �                   @D@X�<ݚ�?             "@�       �                   �A@      �?              @������������������������       ����Q��?             @������������������������       �                     @������������������������       �                     �?������������������������       �                      @������������������������       �                     (@                         �?��S�ۿ?0            �R@                      039@     p�?(             P@                         �?P�Lt�<�?             C@                         �?r�q��?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     @@	                          @8�Z$���?             :@
                        �?@�C��2(�?             6@������������������������       �                     &@                         �?"pc�
�?             &@������������������������       �                     �?                         �?z�G�z�?             $@                         :@�<ݚ�?             "@                        �@@      �?             @������������������������       �                      @������������������������       �                      @������������������������       �                     @������������������������       �                     �?                         ;@      �?             @������������������������       �                     �?                      �|�>@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     &@      F                `D�c@�/,Tg�?7             U@      5                   �?�������?.             Q@                       ��S@�㙢�c�?             G@������������������������       �                     &@      "                   9@4�2%ޑ�?            �A@       !                   �?      �?             @������������������������       �                     @������������������������       �                     @#      *                   �?д>��C�?             =@$      )                `f�S@���N8�?             5@%      (                   �?      �?             @&      '                   �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @������������������������       �                     1@+      2                   �?      �?              @,      -                   �?      �?             @������������������������       �                     �?.      1                   �?���Q��?             @/      0                  �H@      �?             @������������������������       �                      @������������������������       �                      @������������������������       �                     �?3      4                  �G@      �?              @������������������������       �                     �?������������������������       �                     �?6      =                   �?�eP*L��?             6@7      8                    @d}h���?
             ,@������������������������       �                      @9      :                   �?�8��8��?	             (@������������������������       �                     "@;      <                  �5@�q�q�?             @������������������������       �                      @������������������������       �                     �?>      E                   �?      �?              @?      @                   �?؇���X�?             @������������������������       �                     �?A      B                `��S@r�q��?             @������������������������       �                     @C      D                �Cj]@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     �?G      H                ���m@      �?	             0@������������������������       �                     $@I      N                   �?r�q��?             @J      K                   �?�q�q�?             @������������������������       �                     �?L      M                �̾w@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @�t�bh�h(h+K ��h-��R�(KMOKK��h[�B�       `z@      r@     0y@      l@      J@     �b@      C@     �`@      A@      W@      2@     �R@      2@     @P@      1@     @P@              @      1@     �M@       @              .@     �M@      (@      K@      &@      D@       @      D@              @       @     �B@       @      3@      �?              @      3@              "@      @      $@      @      $@      @      @      @              @      @       @      @              @       @              �?      @      �?                      @              @      �?                      2@      @              �?      ,@               @      �?      @      �?      �?              @      @      @      @                      @      �?                      "@      0@      2@      *@      1@              @      *@      ,@       @      @      @      @      �?              @      @       @      @              �?       @       @       @                       @      @              �?              @      &@      @      "@      @                      "@       @       @      �?              �?       @               @      �?              @      �?      @                      �?      @      E@             �C@      @      @      �?      @      �?                      @      @              ,@      0@      @      0@      @       @       @               @       @       @                       @       @      ,@      �?      &@              &@      �?              �?      @      �?       @      �?      �?      �?                      �?              �?              �?       @             �u@     �R@      &@      0@              @      &@      $@              "@      &@      �?      @      �?       @              @      �?      @                      �?      @             @u@     �M@     �a@      (@      $@             �`@      (@      "@       @               @      "@             �^@      $@      C@      @      B@      @     �@@      @      @      @      @       @       @       @               @       @               @                      @      =@      �?      *@      �?      $@              @      �?       @      �?      �?              0@              @      �?              �?      @               @             @U@      @      T@      @      H@              @@      @      �?       @               @      �?              ?@      �?      =@               @      �?              �?       @              @             �h@     �G@      @      @      @               @      @       @       @               @      h@     �E@      ?@      0@      @      @       @              �?      @               @      �?      @              @      �?              <@      &@      6@      $@      �?      @      �?                      @      5@      @      0@      @      0@      @      (@      @       @      @      @      �?      @                      �?      @      @      @       @      @       @      @      �?      �?      �?      �?                      @      @              @                      �?      @              @      �?       @      �?              �?       @              @             @d@      ;@      W@      6@      @      @      @      �?      @               @      �?      �?      �?      �?                      �?      �?                      @     @U@      2@     @R@      2@     �Q@      2@     �O@      &@      @      @              @      @      �?      @              �?      �?              �?      �?             �L@      @      ,@             �E@      @      A@       @      3@              .@       @      (@              @       @      �?       @              �?      �?      �?      �?                      �?       @              "@      @      @      @      @       @       @       @       @                       @      �?                       @      @      �?      @               @      �?              �?       @               @      @      @              @      @              @      @      @      @      @       @      @      @                      �?       @              (@             �Q@      @     �M@      @     �B@      �?      @      �?      @                      �?      @@              6@      @      4@       @      &@              "@       @      �?               @       @      @       @       @       @               @       @              @              �?               @       @              �?       @      �?       @                      �?      &@              3@     @P@      2@      I@       @      C@              &@       @      ;@      @      @              @      @              @      8@      �?      4@      �?      @      �?      �?              �?      �?                       @              1@      @      @      @      @              �?      @       @       @       @               @       @              �?              �?      �?      �?                      �?      $@      (@      @      &@       @              �?      &@              "@      �?       @               @      �?              @      �?      @      �?      �?              @      �?      @               @      �?              �?       @              �?              �?      .@              $@      �?      @      �?       @              �?      �?      �?      �?                      �?              @�t�bub�       hhubehhub.